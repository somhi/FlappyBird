library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ccfbc187",
    12 => x"86c0c64e",
    13 => x"49ccfbc1",
    14 => x"48f8e9c1",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c087f603",
    18 => x"0087cdf8",
    19 => x"1e87fc98",
    20 => x"1e721e73",
    21 => x"ca048bc1",
    22 => x"11481287",
    23 => x"8887c402",
    24 => x"2687f102",
    25 => x"264b264a",
    26 => x"48731e4f",
    27 => x"02a97381",
    28 => x"531287c5",
    29 => x"2687f605",
    30 => x"66c41e4f",
    31 => x"1248714a",
    32 => x"87fb0551",
    33 => x"ff1e4f26",
    34 => x"ffc348d4",
    35 => x"c4516878",
    36 => x"88c14866",
    37 => x"7058a6c8",
    38 => x"87eb0598",
    39 => x"731e4f26",
    40 => x"4bd4ff1e",
    41 => x"6b7bffc3",
    42 => x"7bffc34a",
    43 => x"32c8496b",
    44 => x"ffc3b172",
    45 => x"c84a6b7b",
    46 => x"c3b27131",
    47 => x"496b7bff",
    48 => x"b17232c8",
    49 => x"87c44871",
    50 => x"4c264d26",
    51 => x"4f264b26",
    52 => x"5c5b5e0e",
    53 => x"4a710e5d",
    54 => x"724cd4ff",
    55 => x"99ffc349",
    56 => x"e9c17c71",
    57 => x"c805bff8",
    58 => x"4866d087",
    59 => x"a6d430c9",
    60 => x"4966d058",
    61 => x"ffc329d8",
    62 => x"d07c7199",
    63 => x"29d04966",
    64 => x"7199ffc3",
    65 => x"4966d07c",
    66 => x"ffc329c8",
    67 => x"d07c7199",
    68 => x"ffc34966",
    69 => x"727c7199",
    70 => x"c329d049",
    71 => x"7c7199ff",
    72 => x"f0c94b6c",
    73 => x"ffc34dff",
    74 => x"87d005ab",
    75 => x"6c7cffc3",
    76 => x"028dc14b",
    77 => x"ffc387c6",
    78 => x"87f002ab",
    79 => x"c7fe4873",
    80 => x"d4ff1e87",
    81 => x"48d0ff4a",
    82 => x"c378d1c4",
    83 => x"89c17aff",
    84 => x"2687f805",
    85 => x"1e731e4f",
    86 => x"eec54b71",
    87 => x"ff4adfcd",
    88 => x"ffc348d4",
    89 => x"c3486878",
    90 => x"c502a8fe",
    91 => x"058ac187",
    92 => x"9a7287ed",
    93 => x"c087c505",
    94 => x"87eac048",
    95 => x"cc029b73",
    96 => x"1e66c887",
    97 => x"fdfb4973",
    98 => x"c686c487",
    99 => x"4966c887",
   100 => x"ff87eefe",
   101 => x"ffc348d4",
   102 => x"9b737878",
   103 => x"ff87c505",
   104 => x"78d048d0",
   105 => x"e3fc48c1",
   106 => x"1e731e87",
   107 => x"4bc04a71",
   108 => x"c348d4ff",
   109 => x"d0ff78ff",
   110 => x"78c3c448",
   111 => x"c348d4ff",
   112 => x"1e7278ff",
   113 => x"c1f0ffc0",
   114 => x"c3fc49d1",
   115 => x"7086c487",
   116 => x"87cd0598",
   117 => x"cc1ec0c8",
   118 => x"f8fd4966",
   119 => x"7086c487",
   120 => x"48d0ff4b",
   121 => x"487378c2",
   122 => x"0e87e1fb",
   123 => x"5d5c5b5e",
   124 => x"c186f80e",
   125 => x"c048d0f2",
   126 => x"c8eac178",
   127 => x"fe49c01e",
   128 => x"86c487e7",
   129 => x"c5059870",
   130 => x"c948c087",
   131 => x"4dc087c7",
   132 => x"e6da7ec1",
   133 => x"eac149bf",
   134 => x"c8714afe",
   135 => x"87eff84b",
   136 => x"c2059870",
   137 => x"da7ec087",
   138 => x"c149bfe2",
   139 => x"714adaeb",
   140 => x"daf84bc8",
   141 => x"05987087",
   142 => x"7ec087c2",
   143 => x"fdc0026e",
   144 => x"cef1c187",
   145 => x"f2c14dbf",
   146 => x"7ebf9fc6",
   147 => x"ead6c548",
   148 => x"87c705a8",
   149 => x"bfcef1c1",
   150 => x"6e87ce4d",
   151 => x"d5e9ca48",
   152 => x"87c502a8",
   153 => x"ecc748c0",
   154 => x"c8eac187",
   155 => x"fc49751e",
   156 => x"86c487f7",
   157 => x"c5059870",
   158 => x"c748c087",
   159 => x"e2da87d7",
   160 => x"ebc149bf",
   161 => x"c8714ada",
   162 => x"87c3f74b",
   163 => x"c8059870",
   164 => x"d0f2c187",
   165 => x"d878c148",
   166 => x"bfe6da87",
   167 => x"feeac149",
   168 => x"4bc8714a",
   169 => x"7087e8f6",
   170 => x"87c50298",
   171 => x"e4c648c0",
   172 => x"c6f2c187",
   173 => x"c149bf97",
   174 => x"cd05a9d5",
   175 => x"c7f2c187",
   176 => x"c249bf97",
   177 => x"c002a9ea",
   178 => x"48c087c5",
   179 => x"c187c6c6",
   180 => x"bf97c8ea",
   181 => x"e9c3487e",
   182 => x"cec002a8",
   183 => x"c3486e87",
   184 => x"c002a8eb",
   185 => x"48c087c5",
   186 => x"c187eac5",
   187 => x"bf97d3ea",
   188 => x"c0059949",
   189 => x"eac187cc",
   190 => x"49bf97d4",
   191 => x"c002a9c2",
   192 => x"48c087c5",
   193 => x"c187cec5",
   194 => x"bf97d5ea",
   195 => x"ccf2c148",
   196 => x"484c7058",
   197 => x"f2c188c1",
   198 => x"eac158d0",
   199 => x"49bf97d6",
   200 => x"eac18175",
   201 => x"4abf97d7",
   202 => x"a17232c8",
   203 => x"ddf6c17e",
   204 => x"c1786e48",
   205 => x"bf97d8ea",
   206 => x"58a6c848",
   207 => x"bfd0f2c1",
   208 => x"87d3c202",
   209 => x"49bfe2da",
   210 => x"4adaebc1",
   211 => x"f34bc871",
   212 => x"987087fd",
   213 => x"87c5c002",
   214 => x"f8c348c0",
   215 => x"c8f2c187",
   216 => x"f6c14cbf",
   217 => x"eac15cf1",
   218 => x"49bf97ed",
   219 => x"eac131c8",
   220 => x"4abf97ec",
   221 => x"eac149a1",
   222 => x"4abf97ee",
   223 => x"a17232d0",
   224 => x"efeac149",
   225 => x"d84abf97",
   226 => x"49a17232",
   227 => x"c19166c4",
   228 => x"81bfddf6",
   229 => x"59e5f6c1",
   230 => x"97f5eac1",
   231 => x"32c84abf",
   232 => x"97f4eac1",
   233 => x"4aa24bbf",
   234 => x"97f6eac1",
   235 => x"33d04bbf",
   236 => x"c14aa273",
   237 => x"bf97f7ea",
   238 => x"d89bcf4b",
   239 => x"4aa27333",
   240 => x"5ae9f6c1",
   241 => x"bfe5f6c1",
   242 => x"748ac24a",
   243 => x"e9f6c192",
   244 => x"78a17248",
   245 => x"c187cac1",
   246 => x"bf97daea",
   247 => x"c131c849",
   248 => x"bf97d9ea",
   249 => x"c149a14a",
   250 => x"c159d8f2",
   251 => x"49bfd4f2",
   252 => x"ffc731c5",
   253 => x"c129c981",
   254 => x"c159f1f6",
   255 => x"bf97dfea",
   256 => x"c132c84a",
   257 => x"bf97deea",
   258 => x"c44aa24b",
   259 => x"826e9266",
   260 => x"5aedf6c1",
   261 => x"48e5f6c1",
   262 => x"f6c178c0",
   263 => x"a17248e1",
   264 => x"f1f6c178",
   265 => x"e5f6c148",
   266 => x"f6c178bf",
   267 => x"f6c148f5",
   268 => x"c178bfe9",
   269 => x"02bfd0f2",
   270 => x"7487c9c0",
   271 => x"7030c448",
   272 => x"87c9c07e",
   273 => x"bfedf6c1",
   274 => x"7030c448",
   275 => x"d4f2c17e",
   276 => x"c1786e48",
   277 => x"268ef848",
   278 => x"264c264d",
   279 => x"0e4f264b",
   280 => x"5d5c5b5e",
   281 => x"c14a710e",
   282 => x"02bfd0f2",
   283 => x"4b7287cb",
   284 => x"4c722bc7",
   285 => x"c99cffc1",
   286 => x"c84b7287",
   287 => x"c34c722b",
   288 => x"f6c19cff",
   289 => x"da83bfdd",
   290 => x"02abbfde",
   291 => x"e2da87d8",
   292 => x"c8eac15b",
   293 => x"f449731e",
   294 => x"86c487cf",
   295 => x"c5059870",
   296 => x"c048c087",
   297 => x"f2c187e6",
   298 => x"d202bfd0",
   299 => x"c4497487",
   300 => x"c8eac191",
   301 => x"cf4d6981",
   302 => x"ffffffff",
   303 => x"7487cb9d",
   304 => x"c191c249",
   305 => x"9f81c8ea",
   306 => x"48754d69",
   307 => x"0e87c8fe",
   308 => x"5d5c5b5e",
   309 => x"7186f40e",
   310 => x"727ec04a",
   311 => x"87d8029a",
   312 => x"48c4eac1",
   313 => x"e9c178c0",
   314 => x"f6c148fc",
   315 => x"c178bff5",
   316 => x"c148c0ea",
   317 => x"78bff1f6",
   318 => x"48e5f2c1",
   319 => x"f2c150c0",
   320 => x"c149bfd4",
   321 => x"4abfc4ea",
   322 => x"c303aa71",
   323 => x"497287f8",
   324 => x"df0599cf",
   325 => x"c8eac187",
   326 => x"fce9c11e",
   327 => x"e9c149bf",
   328 => x"a1c148fc",
   329 => x"c0f27178",
   330 => x"da86c487",
   331 => x"eac148da",
   332 => x"87ca78c8",
   333 => x"48bfdada",
   334 => x"da80e0c0",
   335 => x"eac158de",
   336 => x"c148bfc4",
   337 => x"c8eac180",
   338 => x"069a2758",
   339 => x"97bf0000",
   340 => x"029d4dbf",
   341 => x"c387dfc2",
   342 => x"c202ade5",
   343 => x"dada87d8",
   344 => x"a3cb4bbf",
   345 => x"cf4c1149",
   346 => x"d2c105ac",
   347 => x"df497587",
   348 => x"cd89c199",
   349 => x"d8f2c191",
   350 => x"4aa3c181",
   351 => x"a3c35112",
   352 => x"c551124a",
   353 => x"51124aa3",
   354 => x"124aa3c7",
   355 => x"4aa3c951",
   356 => x"a3ce5112",
   357 => x"d051124a",
   358 => x"51124aa3",
   359 => x"124aa3d2",
   360 => x"4aa3d451",
   361 => x"a3d65112",
   362 => x"d851124a",
   363 => x"51124aa3",
   364 => x"124aa3dc",
   365 => x"4aa3de51",
   366 => x"7ec15112",
   367 => x"7487f7c0",
   368 => x"0599c849",
   369 => x"7487e8c0",
   370 => x"0599d049",
   371 => x"66dc87cf",
   372 => x"7387ca02",
   373 => x"0f66dc49",
   374 => x"d2029870",
   375 => x"c0056e87",
   376 => x"f2c187c6",
   377 => x"50c048d8",
   378 => x"48bfdada",
   379 => x"c187e6c2",
   380 => x"c048e5f2",
   381 => x"f2c17e50",
   382 => x"c149bfd4",
   383 => x"4abfc4ea",
   384 => x"fc04aa71",
   385 => x"f6c187c8",
   386 => x"c005bff5",
   387 => x"f2c187c8",
   388 => x"c102bfd0",
   389 => x"deda87fd",
   390 => x"c178ff48",
   391 => x"49bfc0ea",
   392 => x"7087fcf8",
   393 => x"c4eac149",
   394 => x"48a6c459",
   395 => x"bfc0eac1",
   396 => x"d0f2c178",
   397 => x"d8c002bf",
   398 => x"4966c487",
   399 => x"ffffffcf",
   400 => x"02a999f8",
   401 => x"c087c5c0",
   402 => x"87e1c04d",
   403 => x"dcc04dc1",
   404 => x"4966c487",
   405 => x"99f8ffcf",
   406 => x"c8c002a9",
   407 => x"48a6c887",
   408 => x"c5c078c0",
   409 => x"48a6c887",
   410 => x"66c878c1",
   411 => x"059d754d",
   412 => x"c487e0c0",
   413 => x"89c24966",
   414 => x"bfc8f2c1",
   415 => x"f6c1914a",
   416 => x"c14abfe1",
   417 => x"7248fce9",
   418 => x"eac178a1",
   419 => x"78c048c4",
   420 => x"c087ebf9",
   421 => x"f68ef448",
   422 => x"000087fd",
   423 => x"ffff0000",
   424 => x"06aaffff",
   425 => x"06b30000",
   426 => x"41460000",
   427 => x"20323354",
   428 => x"46002020",
   429 => x"36315441",
   430 => x"00202020",
   431 => x"48d4ff1e",
   432 => x"6878ffc3",
   433 => x"1e4f2648",
   434 => x"c348d4ff",
   435 => x"d0ff78ff",
   436 => x"78e1c848",
   437 => x"d448d4ff",
   438 => x"f9f6c178",
   439 => x"bfd4ff48",
   440 => x"1e4f2650",
   441 => x"c048d0ff",
   442 => x"4f2678e0",
   443 => x"87ccff1e",
   444 => x"02994970",
   445 => x"fbc087c6",
   446 => x"87f105a9",
   447 => x"4f264871",
   448 => x"5c5b5e0e",
   449 => x"c04b710e",
   450 => x"87f0fe4c",
   451 => x"02994970",
   452 => x"c087f9c0",
   453 => x"c002a9ec",
   454 => x"fbc087f2",
   455 => x"ebc002a9",
   456 => x"b766cc87",
   457 => x"87c703ac",
   458 => x"c20266d0",
   459 => x"71537187",
   460 => x"87c20299",
   461 => x"c3fe84c1",
   462 => x"99497087",
   463 => x"c087cd02",
   464 => x"c702a9ec",
   465 => x"a9fbc087",
   466 => x"87d5ff05",
   467 => x"c30266d0",
   468 => x"7b97c087",
   469 => x"05a9ecc0",
   470 => x"4a7487c4",
   471 => x"4a7487c5",
   472 => x"728a0ac0",
   473 => x"2687c248",
   474 => x"264c264d",
   475 => x"1e4f264b",
   476 => x"7087c9fd",
   477 => x"b7f0c049",
   478 => x"87ca04a9",
   479 => x"a9b7f9c0",
   480 => x"c087c301",
   481 => x"c1c189f0",
   482 => x"ca04a9b7",
   483 => x"b7dac187",
   484 => x"87c301a9",
   485 => x"7189f7c0",
   486 => x"0e4f2648",
   487 => x"5d5c5b5e",
   488 => x"7186f80e",
   489 => x"fc7ec04c",
   490 => x"4bc087dd",
   491 => x"97c8e1c0",
   492 => x"a9c049bf",
   493 => x"fc87cf04",
   494 => x"83c187f2",
   495 => x"97c8e1c0",
   496 => x"06ab49bf",
   497 => x"e1c087f1",
   498 => x"02bf97c8",
   499 => x"ebfb87cf",
   500 => x"99497087",
   501 => x"c087c602",
   502 => x"f105a9ec",
   503 => x"fb4bc087",
   504 => x"4d7087da",
   505 => x"c887d5fb",
   506 => x"cffb58a6",
   507 => x"c14a7087",
   508 => x"49a4c883",
   509 => x"ad496997",
   510 => x"c087c702",
   511 => x"c005adff",
   512 => x"a4c987e7",
   513 => x"49699749",
   514 => x"02a966c4",
   515 => x"c04887c7",
   516 => x"d405a8ff",
   517 => x"49a4ca87",
   518 => x"aa496997",
   519 => x"c087c602",
   520 => x"c405aaff",
   521 => x"d07ec187",
   522 => x"adecc087",
   523 => x"c087c602",
   524 => x"c405adfb",
   525 => x"c14bc087",
   526 => x"fe026e7e",
   527 => x"e2fa87e1",
   528 => x"f8487387",
   529 => x"87dffc8e",
   530 => x"5b5e0e00",
   531 => x"1e0e5d5c",
   532 => x"4cc04b71",
   533 => x"c004ab4d",
   534 => x"dbde87e7",
   535 => x"029d751e",
   536 => x"4ac087c4",
   537 => x"4ac187c2",
   538 => x"e2f14972",
   539 => x"7086c487",
   540 => x"6e84c17e",
   541 => x"7387c205",
   542 => x"7385c14c",
   543 => x"d9ff06ac",
   544 => x"26486e87",
   545 => x"4c264d26",
   546 => x"4f264b26",
   547 => x"1e4f261e",
   548 => x"4f2648c0",
   549 => x"494a711e",
   550 => x"f9c091cb",
   551 => x"81c881fc",
   552 => x"f6c14811",
   553 => x"f6c158fe",
   554 => x"78c048fe",
   555 => x"d3d549c1",
   556 => x"1e4f2687",
   557 => x"f9c049c0",
   558 => x"4f2687e2",
   559 => x"0299711e",
   560 => x"fbc087d2",
   561 => x"50c048d1",
   562 => x"e2c080f7",
   563 => x"f9c040d4",
   564 => x"87ce78f5",
   565 => x"48cdfbc0",
   566 => x"78eef9c0",
   567 => x"e2c080fc",
   568 => x"4f2678f3",
   569 => x"5c5b5e0e",
   570 => x"4a4c710e",
   571 => x"f9c092cb",
   572 => x"a2c882fc",
   573 => x"4ba2c949",
   574 => x"1e4b6b97",
   575 => x"1e496997",
   576 => x"491282ca",
   577 => x"87dde4c0",
   578 => x"f7d349c0",
   579 => x"c0497487",
   580 => x"f887e4f6",
   581 => x"87eefd8e",
   582 => x"711e731e",
   583 => x"c3ff494b",
   584 => x"fe497387",
   585 => x"49c087fe",
   586 => x"87f0f7c0",
   587 => x"1e87d9fd",
   588 => x"4b711e73",
   589 => x"024aa3c6",
   590 => x"8ac187db",
   591 => x"8a87d602",
   592 => x"87dac102",
   593 => x"fcc0028a",
   594 => x"c0028a87",
   595 => x"028a87e1",
   596 => x"dbc187cb",
   597 => x"fc49c787",
   598 => x"dec187fa",
   599 => x"fef6c187",
   600 => x"cbc102bf",
   601 => x"88c14887",
   602 => x"58c2f7c1",
   603 => x"c187c1c1",
   604 => x"02bfc2f7",
   605 => x"c187f9c0",
   606 => x"48bffef6",
   607 => x"f7c180c1",
   608 => x"ebc058c2",
   609 => x"fef6c187",
   610 => x"89c649bf",
   611 => x"59c2f7c1",
   612 => x"03a9b7c0",
   613 => x"f6c187da",
   614 => x"78c048fe",
   615 => x"f7c187d2",
   616 => x"cb02bfc2",
   617 => x"fef6c187",
   618 => x"80c648bf",
   619 => x"58c2f7c1",
   620 => x"cfd149c0",
   621 => x"c0497387",
   622 => x"fb87fcf3",
   623 => x"5e0e87ca",
   624 => x"710e5c5b",
   625 => x"1e66cc4c",
   626 => x"93cb4b74",
   627 => x"83fcf9c0",
   628 => x"6a4aa3c4",
   629 => x"e0daff49",
   630 => x"cce2c087",
   631 => x"49a3c87b",
   632 => x"c95166d4",
   633 => x"66d849a3",
   634 => x"49a3ca51",
   635 => x"265166dc",
   636 => x"0e87d3fa",
   637 => x"5d5c5b5e",
   638 => x"86d0ff0e",
   639 => x"c459a6d8",
   640 => x"78c048a6",
   641 => x"c4c180c4",
   642 => x"80c47866",
   643 => x"80c478c1",
   644 => x"f7c178c1",
   645 => x"78c148c2",
   646 => x"bffaf6c1",
   647 => x"05a8de48",
   648 => x"eaf987cb",
   649 => x"c8497087",
   650 => x"e0ce59a6",
   651 => x"87d7f287",
   652 => x"f287f9f2",
   653 => x"4c7087c6",
   654 => x"02acfbc0",
   655 => x"d487d0c1",
   656 => x"c2c10566",
   657 => x"1e1ec087",
   658 => x"fbc01ec1",
   659 => x"49c01edf",
   660 => x"c187ebfd",
   661 => x"c44a66d0",
   662 => x"c7496a82",
   663 => x"c1517481",
   664 => x"6a1ed81e",
   665 => x"f281c849",
   666 => x"86d887d6",
   667 => x"4866c4c1",
   668 => x"c701a8c0",
   669 => x"48a6c487",
   670 => x"87ce78c1",
   671 => x"4866c4c1",
   672 => x"a6cc88c1",
   673 => x"f187c358",
   674 => x"a6cc87e2",
   675 => x"7478c248",
   676 => x"f5cc029c",
   677 => x"4866c487",
   678 => x"a866c8c1",
   679 => x"87eacc03",
   680 => x"c048a6d8",
   681 => x"c080c478",
   682 => x"87d0f078",
   683 => x"d0c14c70",
   684 => x"d7c205ac",
   685 => x"7e66dc87",
   686 => x"7087f4f2",
   687 => x"a6e0c049",
   688 => x"87f8ef59",
   689 => x"ecc04c70",
   690 => x"eac105ac",
   691 => x"4966c487",
   692 => x"c0c191cb",
   693 => x"a1c48166",
   694 => x"c84d6a4a",
   695 => x"66dc4aa1",
   696 => x"d4e2c052",
   697 => x"87d4ef79",
   698 => x"029c4c70",
   699 => x"fbc087d8",
   700 => x"87d202ac",
   701 => x"c3ef5574",
   702 => x"9c4c7087",
   703 => x"c087c702",
   704 => x"ff05acfb",
   705 => x"e0c087ee",
   706 => x"55c1c255",
   707 => x"d47d97c0",
   708 => x"a96e4966",
   709 => x"c487db05",
   710 => x"66c84866",
   711 => x"87ca04a8",
   712 => x"c14866c4",
   713 => x"58a6c880",
   714 => x"66c887c8",
   715 => x"cc88c148",
   716 => x"c7ee58a6",
   717 => x"c14c7087",
   718 => x"c805acd0",
   719 => x"4866d087",
   720 => x"a6d480c1",
   721 => x"acd0c158",
   722 => x"87e9fd02",
   723 => x"48a6e0c0",
   724 => x"dc7866d4",
   725 => x"e0c04866",
   726 => x"c805a866",
   727 => x"e4c087ff",
   728 => x"78c048a6",
   729 => x"c048747e",
   730 => x"ecc088fb",
   731 => x"987058a6",
   732 => x"87c4c802",
   733 => x"c088cb48",
   734 => x"7058a6ec",
   735 => x"d0c10298",
   736 => x"88c94887",
   737 => x"58a6ecc0",
   738 => x"c3029870",
   739 => x"c44887d6",
   740 => x"a6ecc088",
   741 => x"02987058",
   742 => x"c14887d0",
   743 => x"a6ecc088",
   744 => x"02987058",
   745 => x"c787fdc2",
   746 => x"a6d887c9",
   747 => x"78f0c048",
   748 => x"7087c9ec",
   749 => x"acecc04c",
   750 => x"87c3c002",
   751 => x"c05ca6dc",
   752 => x"cc02acec",
   753 => x"87f4eb87",
   754 => x"ecc04c70",
   755 => x"f4ff05ac",
   756 => x"acecc087",
   757 => x"87c3c002",
   758 => x"d887e1eb",
   759 => x"66d41e66",
   760 => x"66d41e49",
   761 => x"fbc01e49",
   762 => x"66d41edf",
   763 => x"87cef749",
   764 => x"1eca1ec0",
   765 => x"cb4966dc",
   766 => x"66d8c191",
   767 => x"48a6d881",
   768 => x"d878a1c4",
   769 => x"eb49bf66",
   770 => x"86d887f6",
   771 => x"06a8b7c0",
   772 => x"c187c4c1",
   773 => x"c81ede1e",
   774 => x"eb49bf66",
   775 => x"86c887e2",
   776 => x"c0484970",
   777 => x"a6dc8808",
   778 => x"a8b7c058",
   779 => x"87e7c006",
   780 => x"dd4866d8",
   781 => x"de03a8b7",
   782 => x"49bf6e87",
   783 => x"c08166d8",
   784 => x"66d851e0",
   785 => x"6e81c149",
   786 => x"c1c281bf",
   787 => x"4966d851",
   788 => x"bf6e81c2",
   789 => x"cc51c081",
   790 => x"80c14866",
   791 => x"c158a6d0",
   792 => x"87d4c47e",
   793 => x"dc87c8ec",
   794 => x"c2ec58a6",
   795 => x"a6ecc087",
   796 => x"a8ecc058",
   797 => x"87cac005",
   798 => x"48a6e8c0",
   799 => x"c07866d8",
   800 => x"f7e887c3",
   801 => x"4966c487",
   802 => x"c0c191cb",
   803 => x"80714866",
   804 => x"4a6e7e70",
   805 => x"496e82c8",
   806 => x"66d881ca",
   807 => x"66e8c051",
   808 => x"d881c149",
   809 => x"48c18966",
   810 => x"49703071",
   811 => x"977189c1",
   812 => x"e2fac17a",
   813 => x"66d849bf",
   814 => x"4a6a9729",
   815 => x"c0987148",
   816 => x"6e58a6f0",
   817 => x"6981c449",
   818 => x"66e0c04d",
   819 => x"a866dc48",
   820 => x"87c8c002",
   821 => x"c048a6d8",
   822 => x"87c5c078",
   823 => x"c148a6d8",
   824 => x"1e66d878",
   825 => x"751ee0c0",
   826 => x"87d4e849",
   827 => x"4c7086c8",
   828 => x"06acb7c0",
   829 => x"7487d3c1",
   830 => x"49e0c085",
   831 => x"4b758974",
   832 => x"4ac1f8c0",
   833 => x"e0cdff71",
   834 => x"c085c287",
   835 => x"c14866e4",
   836 => x"a6e8c080",
   837 => x"66ecc058",
   838 => x"7081c149",
   839 => x"c8c002a9",
   840 => x"48a6d887",
   841 => x"c5c078c0",
   842 => x"48a6d887",
   843 => x"66d878c1",
   844 => x"49a4c21e",
   845 => x"7148e0c0",
   846 => x"1e497088",
   847 => x"ffe64975",
   848 => x"c086c887",
   849 => x"ff01a8b7",
   850 => x"e4c087c1",
   851 => x"d1c00266",
   852 => x"c9496e87",
   853 => x"66e4c081",
   854 => x"c0486e51",
   855 => x"c078e4e3",
   856 => x"496e87cc",
   857 => x"51c281c9",
   858 => x"e4c0486e",
   859 => x"7ec178d8",
   860 => x"e587c5c0",
   861 => x"4c7087f6",
   862 => x"f4c0026e",
   863 => x"4866c487",
   864 => x"04a866c8",
   865 => x"c487cbc0",
   866 => x"80c14866",
   867 => x"c058a6c8",
   868 => x"66c887df",
   869 => x"cc88c148",
   870 => x"d4c058a6",
   871 => x"acc6c187",
   872 => x"87c8c005",
   873 => x"c14866cc",
   874 => x"58a6d080",
   875 => x"7087fde4",
   876 => x"4866d04c",
   877 => x"a6d480c1",
   878 => x"029c7458",
   879 => x"c487cbc0",
   880 => x"c8c14866",
   881 => x"f304a866",
   882 => x"d6e487d6",
   883 => x"4866c487",
   884 => x"c003a8c7",
   885 => x"f7c187e5",
   886 => x"78c048c2",
   887 => x"cb4966c4",
   888 => x"66c0c191",
   889 => x"4aa1c481",
   890 => x"52c04a6a",
   891 => x"4866c479",
   892 => x"a6c880c1",
   893 => x"04a8c758",
   894 => x"ff87dbff",
   895 => x"c3ea8ed0",
   896 => x"00203a87",
   897 => x"711e731e",
   898 => x"c6029b4b",
   899 => x"fef6c187",
   900 => x"c778c048",
   901 => x"fef6c11e",
   902 => x"c01e49bf",
   903 => x"c11efcf9",
   904 => x"49bffaf6",
   905 => x"cc87ccef",
   906 => x"faf6c186",
   907 => x"cbea49bf",
   908 => x"029b7387",
   909 => x"f9c087c8",
   910 => x"e3c049fc",
   911 => x"c7e987cb",
   912 => x"f9c51e87",
   913 => x"fe49c187",
   914 => x"f0c287fa",
   915 => x"1e4f2687",
   916 => x"87d1e7c0",
   917 => x"4f2687fa",
   918 => x"fef6c11e",
   919 => x"c178c048",
   920 => x"c048faf6",
   921 => x"87d9ff78",
   922 => x"48c087e5",
   923 => x"20804f26",
   924 => x"74697845",
   925 => x"42208000",
   926 => x"006b6361",
   927 => x"00000894",
   928 => x"00001dc6",
   929 => x"94000000",
   930 => x"e4000008",
   931 => x"0000001d",
   932 => x"08940000",
   933 => x"1e020000",
   934 => x"00000000",
   935 => x"00089400",
   936 => x"001e2000",
   937 => x"00000000",
   938 => x"00000894",
   939 => x"00001e3e",
   940 => x"94000000",
   941 => x"5c000008",
   942 => x"0000001e",
   943 => x"08940000",
   944 => x"1e7a0000",
   945 => x"00000000",
   946 => x"00089400",
   947 => x"00000000",
   948 => x"00000000",
   949 => x"0000092f",
   950 => x"00000000",
   951 => x"4c000000",
   952 => x"2064616f",
   953 => x"1e002e2a",
   954 => x"c048f0fe",
   955 => x"7909cd78",
   956 => x"1e4f2609",
   957 => x"bff0fe1e",
   958 => x"2626487e",
   959 => x"f0fe1e4f",
   960 => x"2678c148",
   961 => x"f0fe1e4f",
   962 => x"2678c048",
   963 => x"4a711e4f",
   964 => x"265252c0",
   965 => x"5b5e0e4f",
   966 => x"f40e5d5c",
   967 => x"974d7186",
   968 => x"a5c17e6d",
   969 => x"486c974c",
   970 => x"6e58a6c8",
   971 => x"a866c448",
   972 => x"ff87c505",
   973 => x"87e6c048",
   974 => x"c287caff",
   975 => x"6c9749a5",
   976 => x"4ba3714b",
   977 => x"974b6b97",
   978 => x"486e7e6c",
   979 => x"a6c880c1",
   980 => x"cc98c758",
   981 => x"977058a6",
   982 => x"87e1fe7c",
   983 => x"8ef44873",
   984 => x"4c264d26",
   985 => x"4f264b26",
   986 => x"5c5b5e0e",
   987 => x"7186f40e",
   988 => x"4a66d84c",
   989 => x"c29affc3",
   990 => x"6c974ba4",
   991 => x"49a17349",
   992 => x"6c975172",
   993 => x"c1486e7e",
   994 => x"58a6c880",
   995 => x"a6cc98c7",
   996 => x"f4547058",
   997 => x"87caff8e",
   998 => x"e8fd1e1e",
   999 => x"4abfe087",
  1000 => x"c0e0c049",
  1001 => x"87cb0299",
  1002 => x"fac11e72",
  1003 => x"f7fe49d8",
  1004 => x"fc86c487",
  1005 => x"7e7087fd",
  1006 => x"2687c2fd",
  1007 => x"c11e4f26",
  1008 => x"fd49d8fa",
  1009 => x"fec087c7",
  1010 => x"dafc49d8",
  1011 => x"87d9c587",
  1012 => x"5e0e4f26",
  1013 => x"0e5d5c5b",
  1014 => x"bff7fac1",
  1015 => x"e6c0c14a",
  1016 => x"724c49bf",
  1017 => x"fc4d71bc",
  1018 => x"4bc087db",
  1019 => x"99d04974",
  1020 => x"7587d502",
  1021 => x"7199d049",
  1022 => x"c11ec01e",
  1023 => x"734af8c6",
  1024 => x"c0491282",
  1025 => x"86c887e4",
  1026 => x"832d2cc1",
  1027 => x"ff04abc8",
  1028 => x"e8fb87da",
  1029 => x"e6c0c187",
  1030 => x"f7fac148",
  1031 => x"4d2678bf",
  1032 => x"4b264c26",
  1033 => x"00004f26",
  1034 => x"ff1e0000",
  1035 => x"e1c848d0",
  1036 => x"48d4ff78",
  1037 => x"66c478c5",
  1038 => x"c387c302",
  1039 => x"66c878e0",
  1040 => x"ff87c602",
  1041 => x"f0c348d4",
  1042 => x"48d4ff78",
  1043 => x"d0ff7871",
  1044 => x"78e1c848",
  1045 => x"2678e0c0",
  1046 => x"5b5e0e4f",
  1047 => x"4c710e5c",
  1048 => x"49d8fac1",
  1049 => x"7087eefa",
  1050 => x"aab7c04a",
  1051 => x"87e3c204",
  1052 => x"05aae0c3",
  1053 => x"c4c187c9",
  1054 => x"78c148dc",
  1055 => x"c387d4c2",
  1056 => x"c905aaf0",
  1057 => x"d8c4c187",
  1058 => x"c178c148",
  1059 => x"c4c187f5",
  1060 => x"c702bfdc",
  1061 => x"c24b7287",
  1062 => x"87c2b3c0",
  1063 => x"9c744b72",
  1064 => x"c187d105",
  1065 => x"1ebfd8c4",
  1066 => x"bfdcc4c1",
  1067 => x"fd49721e",
  1068 => x"86c887f8",
  1069 => x"bfd8c4c1",
  1070 => x"87e0c002",
  1071 => x"b7c44973",
  1072 => x"c5c19129",
  1073 => x"4a7381f8",
  1074 => x"92c29acf",
  1075 => x"307248c1",
  1076 => x"baff4a70",
  1077 => x"98694872",
  1078 => x"87db7970",
  1079 => x"b7c44973",
  1080 => x"c5c19129",
  1081 => x"4a7381f8",
  1082 => x"92c29acf",
  1083 => x"307248c3",
  1084 => x"69484a70",
  1085 => x"c17970b0",
  1086 => x"c048dcc4",
  1087 => x"d8c4c178",
  1088 => x"c178c048",
  1089 => x"f849d8fa",
  1090 => x"4a7087cb",
  1091 => x"03aab7c0",
  1092 => x"c087ddfd",
  1093 => x"87c8fc48",
  1094 => x"00000000",
  1095 => x"00000000",
  1096 => x"494a711e",
  1097 => x"2687f2fc",
  1098 => x"4ac01e4f",
  1099 => x"91c44972",
  1100 => x"81f8c5c1",
  1101 => x"82c179c0",
  1102 => x"04aab7d0",
  1103 => x"4f2687ee",
  1104 => x"5c5b5e0e",
  1105 => x"4d710e5d",
  1106 => x"7587faf6",
  1107 => x"2ab7c44a",
  1108 => x"f8c5c192",
  1109 => x"cf4c7582",
  1110 => x"6a94c29c",
  1111 => x"2b744b49",
  1112 => x"48c29bc3",
  1113 => x"4c703074",
  1114 => x"4874bcff",
  1115 => x"7a709871",
  1116 => x"7387caf6",
  1117 => x"87e6fa48",
  1118 => x"00000000",
  1119 => x"00000000",
  1120 => x"00000000",
  1121 => x"00000000",
  1122 => x"00000000",
  1123 => x"00000000",
  1124 => x"00000000",
  1125 => x"00000000",
  1126 => x"00000000",
  1127 => x"00000000",
  1128 => x"00000000",
  1129 => x"00000000",
  1130 => x"00000000",
  1131 => x"00000000",
  1132 => x"00000000",
  1133 => x"00000000",
  1134 => x"25261e16",
  1135 => x"3e3d362e",
  1136 => x"48d0ff1e",
  1137 => x"7178e1c8",
  1138 => x"08d4ff48",
  1139 => x"4866c478",
  1140 => x"7808d4ff",
  1141 => x"711e4f26",
  1142 => x"1e66c44a",
  1143 => x"49a2e0c1",
  1144 => x"c887ddff",
  1145 => x"b7c84966",
  1146 => x"48d4ff29",
  1147 => x"d0ff7871",
  1148 => x"78e0c048",
  1149 => x"1e4f2626",
  1150 => x"c34ad4ff",
  1151 => x"d0ff7aff",
  1152 => x"78e1c848",
  1153 => x"fac17ade",
  1154 => x"497abfe2",
  1155 => x"7028c848",
  1156 => x"d048717a",
  1157 => x"717a7028",
  1158 => x"7028d848",
  1159 => x"48d0ff7a",
  1160 => x"2678e0c0",
  1161 => x"5b5e0e4f",
  1162 => x"710e5d5c",
  1163 => x"e2fac14c",
  1164 => x"744b4dbf",
  1165 => x"9b66d02b",
  1166 => x"66d483c1",
  1167 => x"87c204ab",
  1168 => x"4a744bc0",
  1169 => x"724966d0",
  1170 => x"75b9ff31",
  1171 => x"72487399",
  1172 => x"484a7030",
  1173 => x"fac1b071",
  1174 => x"dafe58e6",
  1175 => x"264d2687",
  1176 => x"264b264c",
  1177 => x"d0ff1e4f",
  1178 => x"78c9c848",
  1179 => x"d4ff4871",
  1180 => x"4f267808",
  1181 => x"494a711e",
  1182 => x"d0ff87eb",
  1183 => x"2678c848",
  1184 => x"1e731e4f",
  1185 => x"fac14b71",
  1186 => x"c302bff2",
  1187 => x"87ebc287",
  1188 => x"c848d0ff",
  1189 => x"497378c9",
  1190 => x"ffb1e0c0",
  1191 => x"787148d4",
  1192 => x"48e6fac1",
  1193 => x"66c878c0",
  1194 => x"c387c502",
  1195 => x"87c249ff",
  1196 => x"fac149c0",
  1197 => x"66cc59ee",
  1198 => x"c587c602",
  1199 => x"c44ad5d5",
  1200 => x"ffffcf87",
  1201 => x"f2fac14a",
  1202 => x"f2fac15a",
  1203 => x"c478c148",
  1204 => x"264d2687",
  1205 => x"264b264c",
  1206 => x"5b5e0e4f",
  1207 => x"710e5d5c",
  1208 => x"eefac14a",
  1209 => x"9a724cbf",
  1210 => x"4987cb02",
  1211 => x"c9c191c8",
  1212 => x"83714bf7",
  1213 => x"cdc187c4",
  1214 => x"4dc04bf7",
  1215 => x"99744913",
  1216 => x"bfeafac1",
  1217 => x"48d4ffb9",
  1218 => x"b7c17871",
  1219 => x"b7c8852c",
  1220 => x"87e804ad",
  1221 => x"bfe6fac1",
  1222 => x"c180c848",
  1223 => x"fe58eafa",
  1224 => x"731e87ef",
  1225 => x"134b711e",
  1226 => x"cb029a4a",
  1227 => x"fe497287",
  1228 => x"4a1387e7",
  1229 => x"87f5059a",
  1230 => x"1e87dafe",
  1231 => x"bfe6fac1",
  1232 => x"e6fac149",
  1233 => x"78a1c148",
  1234 => x"a9b7c0c4",
  1235 => x"ff87db03",
  1236 => x"fac148d4",
  1237 => x"c178bfea",
  1238 => x"49bfe6fa",
  1239 => x"48e6fac1",
  1240 => x"c478a1c1",
  1241 => x"04a9b7c0",
  1242 => x"d0ff87e5",
  1243 => x"c178c848",
  1244 => x"c048f2fa",
  1245 => x"004f2678",
  1246 => x"00000000",
  1247 => x"00000000",
  1248 => x"5f5f0000",
  1249 => x"00000000",
  1250 => x"03000303",
  1251 => x"14000003",
  1252 => x"7f147f7f",
  1253 => x"0000147f",
  1254 => x"6b6b2e24",
  1255 => x"4c00123a",
  1256 => x"6c18366a",
  1257 => x"30003256",
  1258 => x"77594f7e",
  1259 => x"0040683a",
  1260 => x"03070400",
  1261 => x"00000000",
  1262 => x"633e1c00",
  1263 => x"00000041",
  1264 => x"3e634100",
  1265 => x"0800001c",
  1266 => x"1c1c3e2a",
  1267 => x"00082a3e",
  1268 => x"3e3e0808",
  1269 => x"00000808",
  1270 => x"60e08000",
  1271 => x"00000000",
  1272 => x"08080808",
  1273 => x"00000808",
  1274 => x"60600000",
  1275 => x"40000000",
  1276 => x"0c183060",
  1277 => x"00010306",
  1278 => x"4d597f3e",
  1279 => x"00003e7f",
  1280 => x"7f7f0604",
  1281 => x"00000000",
  1282 => x"59716342",
  1283 => x"0000464f",
  1284 => x"49496322",
  1285 => x"1800367f",
  1286 => x"7f13161c",
  1287 => x"0000107f",
  1288 => x"45456727",
  1289 => x"0000397d",
  1290 => x"494b7e3c",
  1291 => x"00003079",
  1292 => x"79710101",
  1293 => x"0000070f",
  1294 => x"49497f36",
  1295 => x"0000367f",
  1296 => x"69494f06",
  1297 => x"00001e3f",
  1298 => x"66660000",
  1299 => x"00000000",
  1300 => x"66e68000",
  1301 => x"00000000",
  1302 => x"14140808",
  1303 => x"00002222",
  1304 => x"14141414",
  1305 => x"00001414",
  1306 => x"14142222",
  1307 => x"00000808",
  1308 => x"59510302",
  1309 => x"3e00060f",
  1310 => x"555d417f",
  1311 => x"00001e1f",
  1312 => x"09097f7e",
  1313 => x"00007e7f",
  1314 => x"49497f7f",
  1315 => x"0000367f",
  1316 => x"41633e1c",
  1317 => x"00004141",
  1318 => x"63417f7f",
  1319 => x"00001c3e",
  1320 => x"49497f7f",
  1321 => x"00004141",
  1322 => x"09097f7f",
  1323 => x"00000101",
  1324 => x"49417f3e",
  1325 => x"00007a7b",
  1326 => x"08087f7f",
  1327 => x"00007f7f",
  1328 => x"7f7f4100",
  1329 => x"00000041",
  1330 => x"40406020",
  1331 => x"7f003f7f",
  1332 => x"361c087f",
  1333 => x"00004163",
  1334 => x"40407f7f",
  1335 => x"7f004040",
  1336 => x"060c067f",
  1337 => x"7f007f7f",
  1338 => x"180c067f",
  1339 => x"00007f7f",
  1340 => x"41417f3e",
  1341 => x"00003e7f",
  1342 => x"09097f7f",
  1343 => x"3e00060f",
  1344 => x"7f61417f",
  1345 => x"0000407e",
  1346 => x"19097f7f",
  1347 => x"0000667f",
  1348 => x"594d6f26",
  1349 => x"0000327b",
  1350 => x"7f7f0101",
  1351 => x"00000101",
  1352 => x"40407f3f",
  1353 => x"00003f7f",
  1354 => x"70703f0f",
  1355 => x"7f000f3f",
  1356 => x"3018307f",
  1357 => x"41007f7f",
  1358 => x"1c1c3663",
  1359 => x"01416336",
  1360 => x"7c7c0603",
  1361 => x"61010306",
  1362 => x"474d5971",
  1363 => x"00004143",
  1364 => x"417f7f00",
  1365 => x"01000041",
  1366 => x"180c0603",
  1367 => x"00406030",
  1368 => x"7f414100",
  1369 => x"0800007f",
  1370 => x"0603060c",
  1371 => x"8000080c",
  1372 => x"80808080",
  1373 => x"00008080",
  1374 => x"07030000",
  1375 => x"00000004",
  1376 => x"54547420",
  1377 => x"0000787c",
  1378 => x"44447f7f",
  1379 => x"0000387c",
  1380 => x"44447c38",
  1381 => x"00000044",
  1382 => x"44447c38",
  1383 => x"00007f7f",
  1384 => x"54547c38",
  1385 => x"0000185c",
  1386 => x"057f7e04",
  1387 => x"00000005",
  1388 => x"a4a4bc18",
  1389 => x"00007cfc",
  1390 => x"04047f7f",
  1391 => x"0000787c",
  1392 => x"7d3d0000",
  1393 => x"00000040",
  1394 => x"fd808080",
  1395 => x"0000007d",
  1396 => x"38107f7f",
  1397 => x"0000446c",
  1398 => x"7f3f0000",
  1399 => x"7c000040",
  1400 => x"0c180c7c",
  1401 => x"0000787c",
  1402 => x"04047c7c",
  1403 => x"0000787c",
  1404 => x"44447c38",
  1405 => x"0000387c",
  1406 => x"2424fcfc",
  1407 => x"0000183c",
  1408 => x"24243c18",
  1409 => x"0000fcfc",
  1410 => x"04047c7c",
  1411 => x"0000080c",
  1412 => x"54545c48",
  1413 => x"00002074",
  1414 => x"447f3f04",
  1415 => x"00000044",
  1416 => x"40407c3c",
  1417 => x"00007c7c",
  1418 => x"60603c1c",
  1419 => x"3c001c3c",
  1420 => x"6030607c",
  1421 => x"44003c7c",
  1422 => x"3810386c",
  1423 => x"0000446c",
  1424 => x"60e0bc1c",
  1425 => x"00001c3c",
  1426 => x"5c746444",
  1427 => x"0000444c",
  1428 => x"773e0808",
  1429 => x"00004141",
  1430 => x"7f7f0000",
  1431 => x"00000000",
  1432 => x"3e774141",
  1433 => x"02000808",
  1434 => x"02030101",
  1435 => x"7f000102",
  1436 => x"7f7f7f7f",
  1437 => x"08007f7f",
  1438 => x"3e1c1c08",
  1439 => x"7f7f7f3e",
  1440 => x"1c3e3e7f",
  1441 => x"0008081c",
  1442 => x"7c7c1810",
  1443 => x"00001018",
  1444 => x"7c7c3010",
  1445 => x"10001030",
  1446 => x"78606030",
  1447 => x"4200061e",
  1448 => x"3c183c66",
  1449 => x"78004266",
  1450 => x"c6c26a38",
  1451 => x"6000386c",
  1452 => x"00600000",
  1453 => x"0e006000",
  1454 => x"5d5c5b5e",
  1455 => x"4c711e0e",
  1456 => x"bfc3fbc1",
  1457 => x"c04bc04d",
  1458 => x"02ab741e",
  1459 => x"a6c487c7",
  1460 => x"c578c048",
  1461 => x"48a6c487",
  1462 => x"66c478c1",
  1463 => x"ee49731e",
  1464 => x"86c887df",
  1465 => x"ef49e0c0",
  1466 => x"a5c487ef",
  1467 => x"f0496a4a",
  1468 => x"c6f187f0",
  1469 => x"c185cb87",
  1470 => x"abb7c883",
  1471 => x"87c7ff04",
  1472 => x"264d2626",
  1473 => x"264b264c",
  1474 => x"4a711e4f",
  1475 => x"5ac7fbc1",
  1476 => x"48c7fbc1",
  1477 => x"fe4978c7",
  1478 => x"4f2687dd",
  1479 => x"711e731e",
  1480 => x"aab7c04a",
  1481 => x"c187d303",
  1482 => x"05bfdbe8",
  1483 => x"4bc187c4",
  1484 => x"4bc087c2",
  1485 => x"5bdfe8c1",
  1486 => x"e8c187c4",
  1487 => x"e8c15adf",
  1488 => x"c14abfdb",
  1489 => x"a2c0c19a",
  1490 => x"87e8ec49",
  1491 => x"e8c148fc",
  1492 => x"fe78bfdb",
  1493 => x"711e87ef",
  1494 => x"1e66c44a",
  1495 => x"f5e94972",
  1496 => x"4f262687",
  1497 => x"dbe8c11e",
  1498 => x"f3e649bf",
  1499 => x"fbfac187",
  1500 => x"78bfe848",
  1501 => x"48f7fac1",
  1502 => x"c178bfec",
  1503 => x"4abffbfa",
  1504 => x"99ffc349",
  1505 => x"722ab7c8",
  1506 => x"c1b07148",
  1507 => x"2658c3fb",
  1508 => x"5b5e0e4f",
  1509 => x"710e5d5c",
  1510 => x"87c8ff4b",
  1511 => x"48f6fac1",
  1512 => x"497350c0",
  1513 => x"7087d9e6",
  1514 => x"9cc24c49",
  1515 => x"c949eecb",
  1516 => x"497087f1",
  1517 => x"f6fac14d",
  1518 => x"c105bf97",
  1519 => x"66d087e2",
  1520 => x"fffac149",
  1521 => x"d60599bf",
  1522 => x"4966d487",
  1523 => x"bff7fac1",
  1524 => x"87cb0599",
  1525 => x"e7e54973",
  1526 => x"02987087",
  1527 => x"c187c1c1",
  1528 => x"87c0fe4c",
  1529 => x"c6c94975",
  1530 => x"02987087",
  1531 => x"fac187c6",
  1532 => x"50c148f6",
  1533 => x"97f6fac1",
  1534 => x"e3c005bf",
  1535 => x"fffac187",
  1536 => x"66d049bf",
  1537 => x"d6ff0599",
  1538 => x"f7fac187",
  1539 => x"66d449bf",
  1540 => x"caff0599",
  1541 => x"e4497387",
  1542 => x"987087e6",
  1543 => x"87fffe05",
  1544 => x"dcfb4874",
  1545 => x"5b5e0e87",
  1546 => x"f40e5d5c",
  1547 => x"4c4dc086",
  1548 => x"c47ebfec",
  1549 => x"fbc148a6",
  1550 => x"c178bfc3",
  1551 => x"c71ec01e",
  1552 => x"87cdfd49",
  1553 => x"987086c8",
  1554 => x"ff87cd02",
  1555 => x"87ccfb49",
  1556 => x"e349dac1",
  1557 => x"4dc187ea",
  1558 => x"97f6fac1",
  1559 => x"87c302bf",
  1560 => x"c187e5c7",
  1561 => x"4bbffbfa",
  1562 => x"bfdbe8c1",
  1563 => x"87e9c005",
  1564 => x"e349fdc3",
  1565 => x"fac387ca",
  1566 => x"87c4e349",
  1567 => x"ffc34973",
  1568 => x"c01e7199",
  1569 => x"87cefb49",
  1570 => x"b7c84973",
  1571 => x"c11e7129",
  1572 => x"87c2fb49",
  1573 => x"f9c586c8",
  1574 => x"fffac187",
  1575 => x"029b4bbf",
  1576 => x"e8c187dd",
  1577 => x"c649bfd7",
  1578 => x"987087c5",
  1579 => x"c087c405",
  1580 => x"c287d24b",
  1581 => x"eac549e0",
  1582 => x"dbe8c187",
  1583 => x"c187c658",
  1584 => x"c048d7e8",
  1585 => x"c2497378",
  1586 => x"87cd0599",
  1587 => x"e149ebc3",
  1588 => x"497087ee",
  1589 => x"c20299c2",
  1590 => x"734cfb87",
  1591 => x"0599c149",
  1592 => x"f4c387cd",
  1593 => x"87d8e149",
  1594 => x"99c24970",
  1595 => x"fa87c202",
  1596 => x"c849734c",
  1597 => x"87cd0599",
  1598 => x"e149f5c3",
  1599 => x"497087c2",
  1600 => x"d40299c2",
  1601 => x"c7fbc187",
  1602 => x"87c902bf",
  1603 => x"c188c148",
  1604 => x"c258cbfb",
  1605 => x"c14cff87",
  1606 => x"c449734d",
  1607 => x"87cd0599",
  1608 => x"e049f2c3",
  1609 => x"497087da",
  1610 => x"db0299c2",
  1611 => x"c7fbc187",
  1612 => x"c7487ebf",
  1613 => x"cb03a8b7",
  1614 => x"c1486e87",
  1615 => x"cbfbc180",
  1616 => x"87c2c058",
  1617 => x"4dc14cfe",
  1618 => x"ff49fdc3",
  1619 => x"7087f1df",
  1620 => x"0299c249",
  1621 => x"fbc187d5",
  1622 => x"c002bfc7",
  1623 => x"fbc187c9",
  1624 => x"78c048c7",
  1625 => x"fd87c2c0",
  1626 => x"c34dc14c",
  1627 => x"dfff49fa",
  1628 => x"497087ce",
  1629 => x"d90299c2",
  1630 => x"c7fbc187",
  1631 => x"b7c748bf",
  1632 => x"c9c003a8",
  1633 => x"c7fbc187",
  1634 => x"c078c748",
  1635 => x"4cfc87c2",
  1636 => x"b7c04dc1",
  1637 => x"d1c003ac",
  1638 => x"4a66c487",
  1639 => x"6a82d8c1",
  1640 => x"87c6c002",
  1641 => x"49744b6a",
  1642 => x"1ec00f73",
  1643 => x"c11ef0c3",
  1644 => x"dcf749da",
  1645 => x"7086c887",
  1646 => x"e2c00298",
  1647 => x"48a6c887",
  1648 => x"bfc7fbc1",
  1649 => x"4966c878",
  1650 => x"66c491cb",
  1651 => x"70807148",
  1652 => x"02bf6e7e",
  1653 => x"6e87c8c0",
  1654 => x"66c84bbf",
  1655 => x"750f7349",
  1656 => x"c8c0029d",
  1657 => x"c7fbc187",
  1658 => x"caf349bf",
  1659 => x"dfe8c187",
  1660 => x"ddc002bf",
  1661 => x"f6c04987",
  1662 => x"02987087",
  1663 => x"c187d3c0",
  1664 => x"49bfc7fb",
  1665 => x"c087f0f2",
  1666 => x"87d0f449",
  1667 => x"48dfe8c1",
  1668 => x"8ef478c0",
  1669 => x"0087eaf3",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"1e000000",
  1673 => x"c8ff4a71",
  1674 => x"a17249bf",
  1675 => x"1e4f2648",
  1676 => x"89bfc8ff",
  1677 => x"c0c0c0fe",
  1678 => x"01a9c0c0",
  1679 => x"4ac087c4",
  1680 => x"4ac187c2",
  1681 => x"4f264872",
  1682 => x"f1e9c11e",
  1683 => x"b9c149bf",
  1684 => x"59f5e9c1",
  1685 => x"c348d4ff",
  1686 => x"d0ff78ff",
  1687 => x"78e1c848",
  1688 => x"c148d4ff",
  1689 => x"7131c478",
  1690 => x"48d0ff78",
  1691 => x"2678e0c0",
  1692 => x"0000004f",
  1693 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
