
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"fb",x"c1",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"cc",x"fb",x"c1"),
    14 => (x"48",x"f8",x"e9",x"c1"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c0",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"cd",x"f8"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"72",x"1e",x"73"),
    21 => (x"ca",x"04",x"8b",x"c1"),
    22 => (x"11",x"48",x"12",x"87"),
    23 => (x"88",x"87",x"c4",x"02"),
    24 => (x"26",x"87",x"f1",x"02"),
    25 => (x"26",x"4b",x"26",x"4a"),
    26 => (x"48",x"73",x"1e",x"4f"),
    27 => (x"02",x"a9",x"73",x"81"),
    28 => (x"53",x"12",x"87",x"c5"),
    29 => (x"26",x"87",x"f6",x"05"),
    30 => (x"66",x"c4",x"1e",x"4f"),
    31 => (x"12",x"48",x"71",x"4a"),
    32 => (x"87",x"fb",x"05",x"51"),
    33 => (x"ff",x"1e",x"4f",x"26"),
    34 => (x"ff",x"c3",x"48",x"d4"),
    35 => (x"c4",x"51",x"68",x"78"),
    36 => (x"88",x"c1",x"48",x"66"),
    37 => (x"70",x"58",x"a6",x"c8"),
    38 => (x"87",x"eb",x"05",x"98"),
    39 => (x"73",x"1e",x"4f",x"26"),
    40 => (x"4b",x"d4",x"ff",x"1e"),
    41 => (x"6b",x"7b",x"ff",x"c3"),
    42 => (x"7b",x"ff",x"c3",x"4a"),
    43 => (x"32",x"c8",x"49",x"6b"),
    44 => (x"ff",x"c3",x"b1",x"72"),
    45 => (x"c8",x"4a",x"6b",x"7b"),
    46 => (x"c3",x"b2",x"71",x"31"),
    47 => (x"49",x"6b",x"7b",x"ff"),
    48 => (x"b1",x"72",x"32",x"c8"),
    49 => (x"87",x"c4",x"48",x"71"),
    50 => (x"4c",x"26",x"4d",x"26"),
    51 => (x"4f",x"26",x"4b",x"26"),
    52 => (x"5c",x"5b",x"5e",x"0e"),
    53 => (x"4a",x"71",x"0e",x"5d"),
    54 => (x"72",x"4c",x"d4",x"ff"),
    55 => (x"99",x"ff",x"c3",x"49"),
    56 => (x"e9",x"c1",x"7c",x"71"),
    57 => (x"c8",x"05",x"bf",x"f8"),
    58 => (x"48",x"66",x"d0",x"87"),
    59 => (x"a6",x"d4",x"30",x"c9"),
    60 => (x"49",x"66",x"d0",x"58"),
    61 => (x"ff",x"c3",x"29",x"d8"),
    62 => (x"d0",x"7c",x"71",x"99"),
    63 => (x"29",x"d0",x"49",x"66"),
    64 => (x"71",x"99",x"ff",x"c3"),
    65 => (x"49",x"66",x"d0",x"7c"),
    66 => (x"ff",x"c3",x"29",x"c8"),
    67 => (x"d0",x"7c",x"71",x"99"),
    68 => (x"ff",x"c3",x"49",x"66"),
    69 => (x"72",x"7c",x"71",x"99"),
    70 => (x"c3",x"29",x"d0",x"49"),
    71 => (x"7c",x"71",x"99",x"ff"),
    72 => (x"f0",x"c9",x"4b",x"6c"),
    73 => (x"ff",x"c3",x"4d",x"ff"),
    74 => (x"87",x"d0",x"05",x"ab"),
    75 => (x"6c",x"7c",x"ff",x"c3"),
    76 => (x"02",x"8d",x"c1",x"4b"),
    77 => (x"ff",x"c3",x"87",x"c6"),
    78 => (x"87",x"f0",x"02",x"ab"),
    79 => (x"c7",x"fe",x"48",x"73"),
    80 => (x"d4",x"ff",x"1e",x"87"),
    81 => (x"48",x"d0",x"ff",x"4a"),
    82 => (x"c3",x"78",x"d1",x"c4"),
    83 => (x"89",x"c1",x"7a",x"ff"),
    84 => (x"26",x"87",x"f8",x"05"),
    85 => (x"1e",x"73",x"1e",x"4f"),
    86 => (x"ee",x"c5",x"4b",x"71"),
    87 => (x"ff",x"4a",x"df",x"cd"),
    88 => (x"ff",x"c3",x"48",x"d4"),
    89 => (x"c3",x"48",x"68",x"78"),
    90 => (x"c5",x"02",x"a8",x"fe"),
    91 => (x"05",x"8a",x"c1",x"87"),
    92 => (x"9a",x"72",x"87",x"ed"),
    93 => (x"c0",x"87",x"c5",x"05"),
    94 => (x"87",x"ea",x"c0",x"48"),
    95 => (x"cc",x"02",x"9b",x"73"),
    96 => (x"1e",x"66",x"c8",x"87"),
    97 => (x"fd",x"fb",x"49",x"73"),
    98 => (x"c6",x"86",x"c4",x"87"),
    99 => (x"49",x"66",x"c8",x"87"),
   100 => (x"ff",x"87",x"ee",x"fe"),
   101 => (x"ff",x"c3",x"48",x"d4"),
   102 => (x"9b",x"73",x"78",x"78"),
   103 => (x"ff",x"87",x"c5",x"05"),
   104 => (x"78",x"d0",x"48",x"d0"),
   105 => (x"e3",x"fc",x"48",x"c1"),
   106 => (x"1e",x"73",x"1e",x"87"),
   107 => (x"4b",x"c0",x"4a",x"71"),
   108 => (x"c3",x"48",x"d4",x"ff"),
   109 => (x"d0",x"ff",x"78",x"ff"),
   110 => (x"78",x"c3",x"c4",x"48"),
   111 => (x"c3",x"48",x"d4",x"ff"),
   112 => (x"1e",x"72",x"78",x"ff"),
   113 => (x"c1",x"f0",x"ff",x"c0"),
   114 => (x"c3",x"fc",x"49",x"d1"),
   115 => (x"70",x"86",x"c4",x"87"),
   116 => (x"87",x"cd",x"05",x"98"),
   117 => (x"cc",x"1e",x"c0",x"c8"),
   118 => (x"f8",x"fd",x"49",x"66"),
   119 => (x"70",x"86",x"c4",x"87"),
   120 => (x"48",x"d0",x"ff",x"4b"),
   121 => (x"48",x"73",x"78",x"c2"),
   122 => (x"0e",x"87",x"e1",x"fb"),
   123 => (x"5d",x"5c",x"5b",x"5e"),
   124 => (x"c1",x"86",x"f8",x"0e"),
   125 => (x"c0",x"48",x"d0",x"f2"),
   126 => (x"c8",x"ea",x"c1",x"78"),
   127 => (x"fe",x"49",x"c0",x"1e"),
   128 => (x"86",x"c4",x"87",x"e7"),
   129 => (x"c5",x"05",x"98",x"70"),
   130 => (x"c9",x"48",x"c0",x"87"),
   131 => (x"4d",x"c0",x"87",x"c7"),
   132 => (x"e6",x"da",x"7e",x"c1"),
   133 => (x"ea",x"c1",x"49",x"bf"),
   134 => (x"c8",x"71",x"4a",x"fe"),
   135 => (x"87",x"ef",x"f8",x"4b"),
   136 => (x"c2",x"05",x"98",x"70"),
   137 => (x"da",x"7e",x"c0",x"87"),
   138 => (x"c1",x"49",x"bf",x"e2"),
   139 => (x"71",x"4a",x"da",x"eb"),
   140 => (x"da",x"f8",x"4b",x"c8"),
   141 => (x"05",x"98",x"70",x"87"),
   142 => (x"7e",x"c0",x"87",x"c2"),
   143 => (x"fd",x"c0",x"02",x"6e"),
   144 => (x"ce",x"f1",x"c1",x"87"),
   145 => (x"f2",x"c1",x"4d",x"bf"),
   146 => (x"7e",x"bf",x"9f",x"c6"),
   147 => (x"ea",x"d6",x"c5",x"48"),
   148 => (x"87",x"c7",x"05",x"a8"),
   149 => (x"bf",x"ce",x"f1",x"c1"),
   150 => (x"6e",x"87",x"ce",x"4d"),
   151 => (x"d5",x"e9",x"ca",x"48"),
   152 => (x"87",x"c5",x"02",x"a8"),
   153 => (x"ec",x"c7",x"48",x"c0"),
   154 => (x"c8",x"ea",x"c1",x"87"),
   155 => (x"fc",x"49",x"75",x"1e"),
   156 => (x"86",x"c4",x"87",x"f7"),
   157 => (x"c5",x"05",x"98",x"70"),
   158 => (x"c7",x"48",x"c0",x"87"),
   159 => (x"e2",x"da",x"87",x"d7"),
   160 => (x"eb",x"c1",x"49",x"bf"),
   161 => (x"c8",x"71",x"4a",x"da"),
   162 => (x"87",x"c3",x"f7",x"4b"),
   163 => (x"c8",x"05",x"98",x"70"),
   164 => (x"d0",x"f2",x"c1",x"87"),
   165 => (x"d8",x"78",x"c1",x"48"),
   166 => (x"bf",x"e6",x"da",x"87"),
   167 => (x"fe",x"ea",x"c1",x"49"),
   168 => (x"4b",x"c8",x"71",x"4a"),
   169 => (x"70",x"87",x"e8",x"f6"),
   170 => (x"87",x"c5",x"02",x"98"),
   171 => (x"e4",x"c6",x"48",x"c0"),
   172 => (x"c6",x"f2",x"c1",x"87"),
   173 => (x"c1",x"49",x"bf",x"97"),
   174 => (x"cd",x"05",x"a9",x"d5"),
   175 => (x"c7",x"f2",x"c1",x"87"),
   176 => (x"c2",x"49",x"bf",x"97"),
   177 => (x"c0",x"02",x"a9",x"ea"),
   178 => (x"48",x"c0",x"87",x"c5"),
   179 => (x"c1",x"87",x"c6",x"c6"),
   180 => (x"bf",x"97",x"c8",x"ea"),
   181 => (x"e9",x"c3",x"48",x"7e"),
   182 => (x"ce",x"c0",x"02",x"a8"),
   183 => (x"c3",x"48",x"6e",x"87"),
   184 => (x"c0",x"02",x"a8",x"eb"),
   185 => (x"48",x"c0",x"87",x"c5"),
   186 => (x"c1",x"87",x"ea",x"c5"),
   187 => (x"bf",x"97",x"d3",x"ea"),
   188 => (x"c0",x"05",x"99",x"49"),
   189 => (x"ea",x"c1",x"87",x"cc"),
   190 => (x"49",x"bf",x"97",x"d4"),
   191 => (x"c0",x"02",x"a9",x"c2"),
   192 => (x"48",x"c0",x"87",x"c5"),
   193 => (x"c1",x"87",x"ce",x"c5"),
   194 => (x"bf",x"97",x"d5",x"ea"),
   195 => (x"cc",x"f2",x"c1",x"48"),
   196 => (x"48",x"4c",x"70",x"58"),
   197 => (x"f2",x"c1",x"88",x"c1"),
   198 => (x"ea",x"c1",x"58",x"d0"),
   199 => (x"49",x"bf",x"97",x"d6"),
   200 => (x"ea",x"c1",x"81",x"75"),
   201 => (x"4a",x"bf",x"97",x"d7"),
   202 => (x"a1",x"72",x"32",x"c8"),
   203 => (x"dd",x"f6",x"c1",x"7e"),
   204 => (x"c1",x"78",x"6e",x"48"),
   205 => (x"bf",x"97",x"d8",x"ea"),
   206 => (x"58",x"a6",x"c8",x"48"),
   207 => (x"bf",x"d0",x"f2",x"c1"),
   208 => (x"87",x"d3",x"c2",x"02"),
   209 => (x"49",x"bf",x"e2",x"da"),
   210 => (x"4a",x"da",x"eb",x"c1"),
   211 => (x"f3",x"4b",x"c8",x"71"),
   212 => (x"98",x"70",x"87",x"fd"),
   213 => (x"87",x"c5",x"c0",x"02"),
   214 => (x"f8",x"c3",x"48",x"c0"),
   215 => (x"c8",x"f2",x"c1",x"87"),
   216 => (x"f6",x"c1",x"4c",x"bf"),
   217 => (x"ea",x"c1",x"5c",x"f1"),
   218 => (x"49",x"bf",x"97",x"ed"),
   219 => (x"ea",x"c1",x"31",x"c8"),
   220 => (x"4a",x"bf",x"97",x"ec"),
   221 => (x"ea",x"c1",x"49",x"a1"),
   222 => (x"4a",x"bf",x"97",x"ee"),
   223 => (x"a1",x"72",x"32",x"d0"),
   224 => (x"ef",x"ea",x"c1",x"49"),
   225 => (x"d8",x"4a",x"bf",x"97"),
   226 => (x"49",x"a1",x"72",x"32"),
   227 => (x"c1",x"91",x"66",x"c4"),
   228 => (x"81",x"bf",x"dd",x"f6"),
   229 => (x"59",x"e5",x"f6",x"c1"),
   230 => (x"97",x"f5",x"ea",x"c1"),
   231 => (x"32",x"c8",x"4a",x"bf"),
   232 => (x"97",x"f4",x"ea",x"c1"),
   233 => (x"4a",x"a2",x"4b",x"bf"),
   234 => (x"97",x"f6",x"ea",x"c1"),
   235 => (x"33",x"d0",x"4b",x"bf"),
   236 => (x"c1",x"4a",x"a2",x"73"),
   237 => (x"bf",x"97",x"f7",x"ea"),
   238 => (x"d8",x"9b",x"cf",x"4b"),
   239 => (x"4a",x"a2",x"73",x"33"),
   240 => (x"5a",x"e9",x"f6",x"c1"),
   241 => (x"bf",x"e5",x"f6",x"c1"),
   242 => (x"74",x"8a",x"c2",x"4a"),
   243 => (x"e9",x"f6",x"c1",x"92"),
   244 => (x"78",x"a1",x"72",x"48"),
   245 => (x"c1",x"87",x"ca",x"c1"),
   246 => (x"bf",x"97",x"da",x"ea"),
   247 => (x"c1",x"31",x"c8",x"49"),
   248 => (x"bf",x"97",x"d9",x"ea"),
   249 => (x"c1",x"49",x"a1",x"4a"),
   250 => (x"c1",x"59",x"d8",x"f2"),
   251 => (x"49",x"bf",x"d4",x"f2"),
   252 => (x"ff",x"c7",x"31",x"c5"),
   253 => (x"c1",x"29",x"c9",x"81"),
   254 => (x"c1",x"59",x"f1",x"f6"),
   255 => (x"bf",x"97",x"df",x"ea"),
   256 => (x"c1",x"32",x"c8",x"4a"),
   257 => (x"bf",x"97",x"de",x"ea"),
   258 => (x"c4",x"4a",x"a2",x"4b"),
   259 => (x"82",x"6e",x"92",x"66"),
   260 => (x"5a",x"ed",x"f6",x"c1"),
   261 => (x"48",x"e5",x"f6",x"c1"),
   262 => (x"f6",x"c1",x"78",x"c0"),
   263 => (x"a1",x"72",x"48",x"e1"),
   264 => (x"f1",x"f6",x"c1",x"78"),
   265 => (x"e5",x"f6",x"c1",x"48"),
   266 => (x"f6",x"c1",x"78",x"bf"),
   267 => (x"f6",x"c1",x"48",x"f5"),
   268 => (x"c1",x"78",x"bf",x"e9"),
   269 => (x"02",x"bf",x"d0",x"f2"),
   270 => (x"74",x"87",x"c9",x"c0"),
   271 => (x"70",x"30",x"c4",x"48"),
   272 => (x"87",x"c9",x"c0",x"7e"),
   273 => (x"bf",x"ed",x"f6",x"c1"),
   274 => (x"70",x"30",x"c4",x"48"),
   275 => (x"d4",x"f2",x"c1",x"7e"),
   276 => (x"c1",x"78",x"6e",x"48"),
   277 => (x"26",x"8e",x"f8",x"48"),
   278 => (x"26",x"4c",x"26",x"4d"),
   279 => (x"0e",x"4f",x"26",x"4b"),
   280 => (x"5d",x"5c",x"5b",x"5e"),
   281 => (x"c1",x"4a",x"71",x"0e"),
   282 => (x"02",x"bf",x"d0",x"f2"),
   283 => (x"4b",x"72",x"87",x"cb"),
   284 => (x"4c",x"72",x"2b",x"c7"),
   285 => (x"c9",x"9c",x"ff",x"c1"),
   286 => (x"c8",x"4b",x"72",x"87"),
   287 => (x"c3",x"4c",x"72",x"2b"),
   288 => (x"f6",x"c1",x"9c",x"ff"),
   289 => (x"da",x"83",x"bf",x"dd"),
   290 => (x"02",x"ab",x"bf",x"de"),
   291 => (x"e2",x"da",x"87",x"d8"),
   292 => (x"c8",x"ea",x"c1",x"5b"),
   293 => (x"f4",x"49",x"73",x"1e"),
   294 => (x"86",x"c4",x"87",x"cf"),
   295 => (x"c5",x"05",x"98",x"70"),
   296 => (x"c0",x"48",x"c0",x"87"),
   297 => (x"f2",x"c1",x"87",x"e6"),
   298 => (x"d2",x"02",x"bf",x"d0"),
   299 => (x"c4",x"49",x"74",x"87"),
   300 => (x"c8",x"ea",x"c1",x"91"),
   301 => (x"cf",x"4d",x"69",x"81"),
   302 => (x"ff",x"ff",x"ff",x"ff"),
   303 => (x"74",x"87",x"cb",x"9d"),
   304 => (x"c1",x"91",x"c2",x"49"),
   305 => (x"9f",x"81",x"c8",x"ea"),
   306 => (x"48",x"75",x"4d",x"69"),
   307 => (x"0e",x"87",x"c8",x"fe"),
   308 => (x"5d",x"5c",x"5b",x"5e"),
   309 => (x"71",x"86",x"f4",x"0e"),
   310 => (x"72",x"7e",x"c0",x"4a"),
   311 => (x"87",x"d8",x"02",x"9a"),
   312 => (x"48",x"c4",x"ea",x"c1"),
   313 => (x"e9",x"c1",x"78",x"c0"),
   314 => (x"f6",x"c1",x"48",x"fc"),
   315 => (x"c1",x"78",x"bf",x"f5"),
   316 => (x"c1",x"48",x"c0",x"ea"),
   317 => (x"78",x"bf",x"f1",x"f6"),
   318 => (x"48",x"e5",x"f2",x"c1"),
   319 => (x"f2",x"c1",x"50",x"c0"),
   320 => (x"c1",x"49",x"bf",x"d4"),
   321 => (x"4a",x"bf",x"c4",x"ea"),
   322 => (x"c3",x"03",x"aa",x"71"),
   323 => (x"49",x"72",x"87",x"f8"),
   324 => (x"df",x"05",x"99",x"cf"),
   325 => (x"c8",x"ea",x"c1",x"87"),
   326 => (x"fc",x"e9",x"c1",x"1e"),
   327 => (x"e9",x"c1",x"49",x"bf"),
   328 => (x"a1",x"c1",x"48",x"fc"),
   329 => (x"c0",x"f2",x"71",x"78"),
   330 => (x"da",x"86",x"c4",x"87"),
   331 => (x"ea",x"c1",x"48",x"da"),
   332 => (x"87",x"ca",x"78",x"c8"),
   333 => (x"48",x"bf",x"da",x"da"),
   334 => (x"da",x"80",x"e0",x"c0"),
   335 => (x"ea",x"c1",x"58",x"de"),
   336 => (x"c1",x"48",x"bf",x"c4"),
   337 => (x"c8",x"ea",x"c1",x"80"),
   338 => (x"06",x"9a",x"27",x"58"),
   339 => (x"97",x"bf",x"00",x"00"),
   340 => (x"02",x"9d",x"4d",x"bf"),
   341 => (x"c3",x"87",x"df",x"c2"),
   342 => (x"c2",x"02",x"ad",x"e5"),
   343 => (x"da",x"da",x"87",x"d8"),
   344 => (x"a3",x"cb",x"4b",x"bf"),
   345 => (x"cf",x"4c",x"11",x"49"),
   346 => (x"d2",x"c1",x"05",x"ac"),
   347 => (x"df",x"49",x"75",x"87"),
   348 => (x"cd",x"89",x"c1",x"99"),
   349 => (x"d8",x"f2",x"c1",x"91"),
   350 => (x"4a",x"a3",x"c1",x"81"),
   351 => (x"a3",x"c3",x"51",x"12"),
   352 => (x"c5",x"51",x"12",x"4a"),
   353 => (x"51",x"12",x"4a",x"a3"),
   354 => (x"12",x"4a",x"a3",x"c7"),
   355 => (x"4a",x"a3",x"c9",x"51"),
   356 => (x"a3",x"ce",x"51",x"12"),
   357 => (x"d0",x"51",x"12",x"4a"),
   358 => (x"51",x"12",x"4a",x"a3"),
   359 => (x"12",x"4a",x"a3",x"d2"),
   360 => (x"4a",x"a3",x"d4",x"51"),
   361 => (x"a3",x"d6",x"51",x"12"),
   362 => (x"d8",x"51",x"12",x"4a"),
   363 => (x"51",x"12",x"4a",x"a3"),
   364 => (x"12",x"4a",x"a3",x"dc"),
   365 => (x"4a",x"a3",x"de",x"51"),
   366 => (x"7e",x"c1",x"51",x"12"),
   367 => (x"74",x"87",x"f7",x"c0"),
   368 => (x"05",x"99",x"c8",x"49"),
   369 => (x"74",x"87",x"e8",x"c0"),
   370 => (x"05",x"99",x"d0",x"49"),
   371 => (x"66",x"dc",x"87",x"cf"),
   372 => (x"73",x"87",x"ca",x"02"),
   373 => (x"0f",x"66",x"dc",x"49"),
   374 => (x"d2",x"02",x"98",x"70"),
   375 => (x"c0",x"05",x"6e",x"87"),
   376 => (x"f2",x"c1",x"87",x"c6"),
   377 => (x"50",x"c0",x"48",x"d8"),
   378 => (x"48",x"bf",x"da",x"da"),
   379 => (x"c1",x"87",x"e6",x"c2"),
   380 => (x"c0",x"48",x"e5",x"f2"),
   381 => (x"f2",x"c1",x"7e",x"50"),
   382 => (x"c1",x"49",x"bf",x"d4"),
   383 => (x"4a",x"bf",x"c4",x"ea"),
   384 => (x"fc",x"04",x"aa",x"71"),
   385 => (x"f6",x"c1",x"87",x"c8"),
   386 => (x"c0",x"05",x"bf",x"f5"),
   387 => (x"f2",x"c1",x"87",x"c8"),
   388 => (x"c1",x"02",x"bf",x"d0"),
   389 => (x"de",x"da",x"87",x"fd"),
   390 => (x"c1",x"78",x"ff",x"48"),
   391 => (x"49",x"bf",x"c0",x"ea"),
   392 => (x"70",x"87",x"fc",x"f8"),
   393 => (x"c4",x"ea",x"c1",x"49"),
   394 => (x"48",x"a6",x"c4",x"59"),
   395 => (x"bf",x"c0",x"ea",x"c1"),
   396 => (x"d0",x"f2",x"c1",x"78"),
   397 => (x"d8",x"c0",x"02",x"bf"),
   398 => (x"49",x"66",x"c4",x"87"),
   399 => (x"ff",x"ff",x"ff",x"cf"),
   400 => (x"02",x"a9",x"99",x"f8"),
   401 => (x"c0",x"87",x"c5",x"c0"),
   402 => (x"87",x"e1",x"c0",x"4d"),
   403 => (x"dc",x"c0",x"4d",x"c1"),
   404 => (x"49",x"66",x"c4",x"87"),
   405 => (x"99",x"f8",x"ff",x"cf"),
   406 => (x"c8",x"c0",x"02",x"a9"),
   407 => (x"48",x"a6",x"c8",x"87"),
   408 => (x"c5",x"c0",x"78",x"c0"),
   409 => (x"48",x"a6",x"c8",x"87"),
   410 => (x"66",x"c8",x"78",x"c1"),
   411 => (x"05",x"9d",x"75",x"4d"),
   412 => (x"c4",x"87",x"e0",x"c0"),
   413 => (x"89",x"c2",x"49",x"66"),
   414 => (x"bf",x"c8",x"f2",x"c1"),
   415 => (x"f6",x"c1",x"91",x"4a"),
   416 => (x"c1",x"4a",x"bf",x"e1"),
   417 => (x"72",x"48",x"fc",x"e9"),
   418 => (x"ea",x"c1",x"78",x"a1"),
   419 => (x"78",x"c0",x"48",x"c4"),
   420 => (x"c0",x"87",x"eb",x"f9"),
   421 => (x"f6",x"8e",x"f4",x"48"),
   422 => (x"00",x"00",x"87",x"fd"),
   423 => (x"ff",x"ff",x"00",x"00"),
   424 => (x"06",x"aa",x"ff",x"ff"),
   425 => (x"06",x"b3",x"00",x"00"),
   426 => (x"41",x"46",x"00",x"00"),
   427 => (x"20",x"32",x"33",x"54"),
   428 => (x"46",x"00",x"20",x"20"),
   429 => (x"36",x"31",x"54",x"41"),
   430 => (x"00",x"20",x"20",x"20"),
   431 => (x"48",x"d4",x"ff",x"1e"),
   432 => (x"68",x"78",x"ff",x"c3"),
   433 => (x"1e",x"4f",x"26",x"48"),
   434 => (x"c3",x"48",x"d4",x"ff"),
   435 => (x"d0",x"ff",x"78",x"ff"),
   436 => (x"78",x"e1",x"c8",x"48"),
   437 => (x"d4",x"48",x"d4",x"ff"),
   438 => (x"f9",x"f6",x"c1",x"78"),
   439 => (x"bf",x"d4",x"ff",x"48"),
   440 => (x"1e",x"4f",x"26",x"50"),
   441 => (x"c0",x"48",x"d0",x"ff"),
   442 => (x"4f",x"26",x"78",x"e0"),
   443 => (x"87",x"cc",x"ff",x"1e"),
   444 => (x"02",x"99",x"49",x"70"),
   445 => (x"fb",x"c0",x"87",x"c6"),
   446 => (x"87",x"f1",x"05",x"a9"),
   447 => (x"4f",x"26",x"48",x"71"),
   448 => (x"5c",x"5b",x"5e",x"0e"),
   449 => (x"c0",x"4b",x"71",x"0e"),
   450 => (x"87",x"f0",x"fe",x"4c"),
   451 => (x"02",x"99",x"49",x"70"),
   452 => (x"c0",x"87",x"f9",x"c0"),
   453 => (x"c0",x"02",x"a9",x"ec"),
   454 => (x"fb",x"c0",x"87",x"f2"),
   455 => (x"eb",x"c0",x"02",x"a9"),
   456 => (x"b7",x"66",x"cc",x"87"),
   457 => (x"87",x"c7",x"03",x"ac"),
   458 => (x"c2",x"02",x"66",x"d0"),
   459 => (x"71",x"53",x"71",x"87"),
   460 => (x"87",x"c2",x"02",x"99"),
   461 => (x"c3",x"fe",x"84",x"c1"),
   462 => (x"99",x"49",x"70",x"87"),
   463 => (x"c0",x"87",x"cd",x"02"),
   464 => (x"c7",x"02",x"a9",x"ec"),
   465 => (x"a9",x"fb",x"c0",x"87"),
   466 => (x"87",x"d5",x"ff",x"05"),
   467 => (x"c3",x"02",x"66",x"d0"),
   468 => (x"7b",x"97",x"c0",x"87"),
   469 => (x"05",x"a9",x"ec",x"c0"),
   470 => (x"4a",x"74",x"87",x"c4"),
   471 => (x"4a",x"74",x"87",x"c5"),
   472 => (x"72",x"8a",x"0a",x"c0"),
   473 => (x"26",x"87",x"c2",x"48"),
   474 => (x"26",x"4c",x"26",x"4d"),
   475 => (x"1e",x"4f",x"26",x"4b"),
   476 => (x"70",x"87",x"c9",x"fd"),
   477 => (x"b7",x"f0",x"c0",x"49"),
   478 => (x"87",x"ca",x"04",x"a9"),
   479 => (x"a9",x"b7",x"f9",x"c0"),
   480 => (x"c0",x"87",x"c3",x"01"),
   481 => (x"c1",x"c1",x"89",x"f0"),
   482 => (x"ca",x"04",x"a9",x"b7"),
   483 => (x"b7",x"da",x"c1",x"87"),
   484 => (x"87",x"c3",x"01",x"a9"),
   485 => (x"71",x"89",x"f7",x"c0"),
   486 => (x"0e",x"4f",x"26",x"48"),
   487 => (x"5d",x"5c",x"5b",x"5e"),
   488 => (x"71",x"86",x"f8",x"0e"),
   489 => (x"fc",x"7e",x"c0",x"4c"),
   490 => (x"4b",x"c0",x"87",x"dd"),
   491 => (x"97",x"c8",x"e1",x"c0"),
   492 => (x"a9",x"c0",x"49",x"bf"),
   493 => (x"fc",x"87",x"cf",x"04"),
   494 => (x"83",x"c1",x"87",x"f2"),
   495 => (x"97",x"c8",x"e1",x"c0"),
   496 => (x"06",x"ab",x"49",x"bf"),
   497 => (x"e1",x"c0",x"87",x"f1"),
   498 => (x"02",x"bf",x"97",x"c8"),
   499 => (x"eb",x"fb",x"87",x"cf"),
   500 => (x"99",x"49",x"70",x"87"),
   501 => (x"c0",x"87",x"c6",x"02"),
   502 => (x"f1",x"05",x"a9",x"ec"),
   503 => (x"fb",x"4b",x"c0",x"87"),
   504 => (x"4d",x"70",x"87",x"da"),
   505 => (x"c8",x"87",x"d5",x"fb"),
   506 => (x"cf",x"fb",x"58",x"a6"),
   507 => (x"c1",x"4a",x"70",x"87"),
   508 => (x"49",x"a4",x"c8",x"83"),
   509 => (x"ad",x"49",x"69",x"97"),
   510 => (x"c0",x"87",x"c7",x"02"),
   511 => (x"c0",x"05",x"ad",x"ff"),
   512 => (x"a4",x"c9",x"87",x"e7"),
   513 => (x"49",x"69",x"97",x"49"),
   514 => (x"02",x"a9",x"66",x"c4"),
   515 => (x"c0",x"48",x"87",x"c7"),
   516 => (x"d4",x"05",x"a8",x"ff"),
   517 => (x"49",x"a4",x"ca",x"87"),
   518 => (x"aa",x"49",x"69",x"97"),
   519 => (x"c0",x"87",x"c6",x"02"),
   520 => (x"c4",x"05",x"aa",x"ff"),
   521 => (x"d0",x"7e",x"c1",x"87"),
   522 => (x"ad",x"ec",x"c0",x"87"),
   523 => (x"c0",x"87",x"c6",x"02"),
   524 => (x"c4",x"05",x"ad",x"fb"),
   525 => (x"c1",x"4b",x"c0",x"87"),
   526 => (x"fe",x"02",x"6e",x"7e"),
   527 => (x"e2",x"fa",x"87",x"e1"),
   528 => (x"f8",x"48",x"73",x"87"),
   529 => (x"87",x"df",x"fc",x"8e"),
   530 => (x"5b",x"5e",x"0e",x"00"),
   531 => (x"1e",x"0e",x"5d",x"5c"),
   532 => (x"4c",x"c0",x"4b",x"71"),
   533 => (x"c0",x"04",x"ab",x"4d"),
   534 => (x"db",x"de",x"87",x"e7"),
   535 => (x"02",x"9d",x"75",x"1e"),
   536 => (x"4a",x"c0",x"87",x"c4"),
   537 => (x"4a",x"c1",x"87",x"c2"),
   538 => (x"e2",x"f1",x"49",x"72"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"6e",x"84",x"c1",x"7e"),
   541 => (x"73",x"87",x"c2",x"05"),
   542 => (x"73",x"85",x"c1",x"4c"),
   543 => (x"d9",x"ff",x"06",x"ac"),
   544 => (x"26",x"48",x"6e",x"87"),
   545 => (x"4c",x"26",x"4d",x"26"),
   546 => (x"4f",x"26",x"4b",x"26"),
   547 => (x"1e",x"4f",x"26",x"1e"),
   548 => (x"4f",x"26",x"48",x"c0"),
   549 => (x"49",x"4a",x"71",x"1e"),
   550 => (x"f9",x"c0",x"91",x"cb"),
   551 => (x"81",x"c8",x"81",x"fc"),
   552 => (x"f6",x"c1",x"48",x"11"),
   553 => (x"f6",x"c1",x"58",x"fe"),
   554 => (x"78",x"c0",x"48",x"fe"),
   555 => (x"d3",x"d5",x"49",x"c1"),
   556 => (x"1e",x"4f",x"26",x"87"),
   557 => (x"f9",x"c0",x"49",x"c0"),
   558 => (x"4f",x"26",x"87",x"e2"),
   559 => (x"02",x"99",x"71",x"1e"),
   560 => (x"fb",x"c0",x"87",x"d2"),
   561 => (x"50",x"c0",x"48",x"d1"),
   562 => (x"e2",x"c0",x"80",x"f7"),
   563 => (x"f9",x"c0",x"40",x"d4"),
   564 => (x"87",x"ce",x"78",x"f5"),
   565 => (x"48",x"cd",x"fb",x"c0"),
   566 => (x"78",x"ee",x"f9",x"c0"),
   567 => (x"e2",x"c0",x"80",x"fc"),
   568 => (x"4f",x"26",x"78",x"f3"),
   569 => (x"5c",x"5b",x"5e",x"0e"),
   570 => (x"4a",x"4c",x"71",x"0e"),
   571 => (x"f9",x"c0",x"92",x"cb"),
   572 => (x"a2",x"c8",x"82",x"fc"),
   573 => (x"4b",x"a2",x"c9",x"49"),
   574 => (x"1e",x"4b",x"6b",x"97"),
   575 => (x"1e",x"49",x"69",x"97"),
   576 => (x"49",x"12",x"82",x"ca"),
   577 => (x"87",x"dd",x"e4",x"c0"),
   578 => (x"f7",x"d3",x"49",x"c0"),
   579 => (x"c0",x"49",x"74",x"87"),
   580 => (x"f8",x"87",x"e4",x"f6"),
   581 => (x"87",x"ee",x"fd",x"8e"),
   582 => (x"71",x"1e",x"73",x"1e"),
   583 => (x"c3",x"ff",x"49",x"4b"),
   584 => (x"fe",x"49",x"73",x"87"),
   585 => (x"49",x"c0",x"87",x"fe"),
   586 => (x"87",x"f0",x"f7",x"c0"),
   587 => (x"1e",x"87",x"d9",x"fd"),
   588 => (x"4b",x"71",x"1e",x"73"),
   589 => (x"02",x"4a",x"a3",x"c6"),
   590 => (x"8a",x"c1",x"87",x"db"),
   591 => (x"8a",x"87",x"d6",x"02"),
   592 => (x"87",x"da",x"c1",x"02"),
   593 => (x"fc",x"c0",x"02",x"8a"),
   594 => (x"c0",x"02",x"8a",x"87"),
   595 => (x"02",x"8a",x"87",x"e1"),
   596 => (x"db",x"c1",x"87",x"cb"),
   597 => (x"fc",x"49",x"c7",x"87"),
   598 => (x"de",x"c1",x"87",x"fa"),
   599 => (x"fe",x"f6",x"c1",x"87"),
   600 => (x"cb",x"c1",x"02",x"bf"),
   601 => (x"88",x"c1",x"48",x"87"),
   602 => (x"58",x"c2",x"f7",x"c1"),
   603 => (x"c1",x"87",x"c1",x"c1"),
   604 => (x"02",x"bf",x"c2",x"f7"),
   605 => (x"c1",x"87",x"f9",x"c0"),
   606 => (x"48",x"bf",x"fe",x"f6"),
   607 => (x"f7",x"c1",x"80",x"c1"),
   608 => (x"eb",x"c0",x"58",x"c2"),
   609 => (x"fe",x"f6",x"c1",x"87"),
   610 => (x"89",x"c6",x"49",x"bf"),
   611 => (x"59",x"c2",x"f7",x"c1"),
   612 => (x"03",x"a9",x"b7",x"c0"),
   613 => (x"f6",x"c1",x"87",x"da"),
   614 => (x"78",x"c0",x"48",x"fe"),
   615 => (x"f7",x"c1",x"87",x"d2"),
   616 => (x"cb",x"02",x"bf",x"c2"),
   617 => (x"fe",x"f6",x"c1",x"87"),
   618 => (x"80",x"c6",x"48",x"bf"),
   619 => (x"58",x"c2",x"f7",x"c1"),
   620 => (x"cf",x"d1",x"49",x"c0"),
   621 => (x"c0",x"49",x"73",x"87"),
   622 => (x"fb",x"87",x"fc",x"f3"),
   623 => (x"5e",x"0e",x"87",x"ca"),
   624 => (x"71",x"0e",x"5c",x"5b"),
   625 => (x"1e",x"66",x"cc",x"4c"),
   626 => (x"93",x"cb",x"4b",x"74"),
   627 => (x"83",x"fc",x"f9",x"c0"),
   628 => (x"6a",x"4a",x"a3",x"c4"),
   629 => (x"e0",x"da",x"ff",x"49"),
   630 => (x"cc",x"e2",x"c0",x"87"),
   631 => (x"49",x"a3",x"c8",x"7b"),
   632 => (x"c9",x"51",x"66",x"d4"),
   633 => (x"66",x"d8",x"49",x"a3"),
   634 => (x"49",x"a3",x"ca",x"51"),
   635 => (x"26",x"51",x"66",x"dc"),
   636 => (x"0e",x"87",x"d3",x"fa"),
   637 => (x"5d",x"5c",x"5b",x"5e"),
   638 => (x"86",x"d0",x"ff",x"0e"),
   639 => (x"c4",x"59",x"a6",x"d8"),
   640 => (x"78",x"c0",x"48",x"a6"),
   641 => (x"c4",x"c1",x"80",x"c4"),
   642 => (x"80",x"c4",x"78",x"66"),
   643 => (x"80",x"c4",x"78",x"c1"),
   644 => (x"f7",x"c1",x"78",x"c1"),
   645 => (x"78",x"c1",x"48",x"c2"),
   646 => (x"bf",x"fa",x"f6",x"c1"),
   647 => (x"05",x"a8",x"de",x"48"),
   648 => (x"ea",x"f9",x"87",x"cb"),
   649 => (x"c8",x"49",x"70",x"87"),
   650 => (x"e0",x"ce",x"59",x"a6"),
   651 => (x"87",x"d7",x"f2",x"87"),
   652 => (x"f2",x"87",x"f9",x"f2"),
   653 => (x"4c",x"70",x"87",x"c6"),
   654 => (x"02",x"ac",x"fb",x"c0"),
   655 => (x"d4",x"87",x"d0",x"c1"),
   656 => (x"c2",x"c1",x"05",x"66"),
   657 => (x"1e",x"1e",x"c0",x"87"),
   658 => (x"fb",x"c0",x"1e",x"c1"),
   659 => (x"49",x"c0",x"1e",x"df"),
   660 => (x"c1",x"87",x"eb",x"fd"),
   661 => (x"c4",x"4a",x"66",x"d0"),
   662 => (x"c7",x"49",x"6a",x"82"),
   663 => (x"c1",x"51",x"74",x"81"),
   664 => (x"6a",x"1e",x"d8",x"1e"),
   665 => (x"f2",x"81",x"c8",x"49"),
   666 => (x"86",x"d8",x"87",x"d6"),
   667 => (x"48",x"66",x"c4",x"c1"),
   668 => (x"c7",x"01",x"a8",x"c0"),
   669 => (x"48",x"a6",x"c4",x"87"),
   670 => (x"87",x"ce",x"78",x"c1"),
   671 => (x"48",x"66",x"c4",x"c1"),
   672 => (x"a6",x"cc",x"88",x"c1"),
   673 => (x"f1",x"87",x"c3",x"58"),
   674 => (x"a6",x"cc",x"87",x"e2"),
   675 => (x"74",x"78",x"c2",x"48"),
   676 => (x"f5",x"cc",x"02",x"9c"),
   677 => (x"48",x"66",x"c4",x"87"),
   678 => (x"a8",x"66",x"c8",x"c1"),
   679 => (x"87",x"ea",x"cc",x"03"),
   680 => (x"c0",x"48",x"a6",x"d8"),
   681 => (x"c0",x"80",x"c4",x"78"),
   682 => (x"87",x"d0",x"f0",x"78"),
   683 => (x"d0",x"c1",x"4c",x"70"),
   684 => (x"d7",x"c2",x"05",x"ac"),
   685 => (x"7e",x"66",x"dc",x"87"),
   686 => (x"70",x"87",x"f4",x"f2"),
   687 => (x"a6",x"e0",x"c0",x"49"),
   688 => (x"87",x"f8",x"ef",x"59"),
   689 => (x"ec",x"c0",x"4c",x"70"),
   690 => (x"ea",x"c1",x"05",x"ac"),
   691 => (x"49",x"66",x"c4",x"87"),
   692 => (x"c0",x"c1",x"91",x"cb"),
   693 => (x"a1",x"c4",x"81",x"66"),
   694 => (x"c8",x"4d",x"6a",x"4a"),
   695 => (x"66",x"dc",x"4a",x"a1"),
   696 => (x"d4",x"e2",x"c0",x"52"),
   697 => (x"87",x"d4",x"ef",x"79"),
   698 => (x"02",x"9c",x"4c",x"70"),
   699 => (x"fb",x"c0",x"87",x"d8"),
   700 => (x"87",x"d2",x"02",x"ac"),
   701 => (x"c3",x"ef",x"55",x"74"),
   702 => (x"9c",x"4c",x"70",x"87"),
   703 => (x"c0",x"87",x"c7",x"02"),
   704 => (x"ff",x"05",x"ac",x"fb"),
   705 => (x"e0",x"c0",x"87",x"ee"),
   706 => (x"55",x"c1",x"c2",x"55"),
   707 => (x"d4",x"7d",x"97",x"c0"),
   708 => (x"a9",x"6e",x"49",x"66"),
   709 => (x"c4",x"87",x"db",x"05"),
   710 => (x"66",x"c8",x"48",x"66"),
   711 => (x"87",x"ca",x"04",x"a8"),
   712 => (x"c1",x"48",x"66",x"c4"),
   713 => (x"58",x"a6",x"c8",x"80"),
   714 => (x"66",x"c8",x"87",x"c8"),
   715 => (x"cc",x"88",x"c1",x"48"),
   716 => (x"c7",x"ee",x"58",x"a6"),
   717 => (x"c1",x"4c",x"70",x"87"),
   718 => (x"c8",x"05",x"ac",x"d0"),
   719 => (x"48",x"66",x"d0",x"87"),
   720 => (x"a6",x"d4",x"80",x"c1"),
   721 => (x"ac",x"d0",x"c1",x"58"),
   722 => (x"87",x"e9",x"fd",x"02"),
   723 => (x"48",x"a6",x"e0",x"c0"),
   724 => (x"dc",x"78",x"66",x"d4"),
   725 => (x"e0",x"c0",x"48",x"66"),
   726 => (x"c8",x"05",x"a8",x"66"),
   727 => (x"e4",x"c0",x"87",x"ff"),
   728 => (x"78",x"c0",x"48",x"a6"),
   729 => (x"c0",x"48",x"74",x"7e"),
   730 => (x"ec",x"c0",x"88",x"fb"),
   731 => (x"98",x"70",x"58",x"a6"),
   732 => (x"87",x"c4",x"c8",x"02"),
   733 => (x"c0",x"88",x"cb",x"48"),
   734 => (x"70",x"58",x"a6",x"ec"),
   735 => (x"d0",x"c1",x"02",x"98"),
   736 => (x"88",x"c9",x"48",x"87"),
   737 => (x"58",x"a6",x"ec",x"c0"),
   738 => (x"c3",x"02",x"98",x"70"),
   739 => (x"c4",x"48",x"87",x"d6"),
   740 => (x"a6",x"ec",x"c0",x"88"),
   741 => (x"02",x"98",x"70",x"58"),
   742 => (x"c1",x"48",x"87",x"d0"),
   743 => (x"a6",x"ec",x"c0",x"88"),
   744 => (x"02",x"98",x"70",x"58"),
   745 => (x"c7",x"87",x"fd",x"c2"),
   746 => (x"a6",x"d8",x"87",x"c9"),
   747 => (x"78",x"f0",x"c0",x"48"),
   748 => (x"70",x"87",x"c9",x"ec"),
   749 => (x"ac",x"ec",x"c0",x"4c"),
   750 => (x"87",x"c3",x"c0",x"02"),
   751 => (x"c0",x"5c",x"a6",x"dc"),
   752 => (x"cc",x"02",x"ac",x"ec"),
   753 => (x"87",x"f4",x"eb",x"87"),
   754 => (x"ec",x"c0",x"4c",x"70"),
   755 => (x"f4",x"ff",x"05",x"ac"),
   756 => (x"ac",x"ec",x"c0",x"87"),
   757 => (x"87",x"c3",x"c0",x"02"),
   758 => (x"d8",x"87",x"e1",x"eb"),
   759 => (x"66",x"d4",x"1e",x"66"),
   760 => (x"66",x"d4",x"1e",x"49"),
   761 => (x"fb",x"c0",x"1e",x"49"),
   762 => (x"66",x"d4",x"1e",x"df"),
   763 => (x"87",x"ce",x"f7",x"49"),
   764 => (x"1e",x"ca",x"1e",x"c0"),
   765 => (x"cb",x"49",x"66",x"dc"),
   766 => (x"66",x"d8",x"c1",x"91"),
   767 => (x"48",x"a6",x"d8",x"81"),
   768 => (x"d8",x"78",x"a1",x"c4"),
   769 => (x"eb",x"49",x"bf",x"66"),
   770 => (x"86",x"d8",x"87",x"f6"),
   771 => (x"06",x"a8",x"b7",x"c0"),
   772 => (x"c1",x"87",x"c4",x"c1"),
   773 => (x"c8",x"1e",x"de",x"1e"),
   774 => (x"eb",x"49",x"bf",x"66"),
   775 => (x"86",x"c8",x"87",x"e2"),
   776 => (x"c0",x"48",x"49",x"70"),
   777 => (x"a6",x"dc",x"88",x"08"),
   778 => (x"a8",x"b7",x"c0",x"58"),
   779 => (x"87",x"e7",x"c0",x"06"),
   780 => (x"dd",x"48",x"66",x"d8"),
   781 => (x"de",x"03",x"a8",x"b7"),
   782 => (x"49",x"bf",x"6e",x"87"),
   783 => (x"c0",x"81",x"66",x"d8"),
   784 => (x"66",x"d8",x"51",x"e0"),
   785 => (x"6e",x"81",x"c1",x"49"),
   786 => (x"c1",x"c2",x"81",x"bf"),
   787 => (x"49",x"66",x"d8",x"51"),
   788 => (x"bf",x"6e",x"81",x"c2"),
   789 => (x"cc",x"51",x"c0",x"81"),
   790 => (x"80",x"c1",x"48",x"66"),
   791 => (x"c1",x"58",x"a6",x"d0"),
   792 => (x"87",x"d4",x"c4",x"7e"),
   793 => (x"dc",x"87",x"c8",x"ec"),
   794 => (x"c2",x"ec",x"58",x"a6"),
   795 => (x"a6",x"ec",x"c0",x"87"),
   796 => (x"a8",x"ec",x"c0",x"58"),
   797 => (x"87",x"ca",x"c0",x"05"),
   798 => (x"48",x"a6",x"e8",x"c0"),
   799 => (x"c0",x"78",x"66",x"d8"),
   800 => (x"f7",x"e8",x"87",x"c3"),
   801 => (x"49",x"66",x"c4",x"87"),
   802 => (x"c0",x"c1",x"91",x"cb"),
   803 => (x"80",x"71",x"48",x"66"),
   804 => (x"4a",x"6e",x"7e",x"70"),
   805 => (x"49",x"6e",x"82",x"c8"),
   806 => (x"66",x"d8",x"81",x"ca"),
   807 => (x"66",x"e8",x"c0",x"51"),
   808 => (x"d8",x"81",x"c1",x"49"),
   809 => (x"48",x"c1",x"89",x"66"),
   810 => (x"49",x"70",x"30",x"71"),
   811 => (x"97",x"71",x"89",x"c1"),
   812 => (x"e2",x"fa",x"c1",x"7a"),
   813 => (x"66",x"d8",x"49",x"bf"),
   814 => (x"4a",x"6a",x"97",x"29"),
   815 => (x"c0",x"98",x"71",x"48"),
   816 => (x"6e",x"58",x"a6",x"f0"),
   817 => (x"69",x"81",x"c4",x"49"),
   818 => (x"66",x"e0",x"c0",x"4d"),
   819 => (x"a8",x"66",x"dc",x"48"),
   820 => (x"87",x"c8",x"c0",x"02"),
   821 => (x"c0",x"48",x"a6",x"d8"),
   822 => (x"87",x"c5",x"c0",x"78"),
   823 => (x"c1",x"48",x"a6",x"d8"),
   824 => (x"1e",x"66",x"d8",x"78"),
   825 => (x"75",x"1e",x"e0",x"c0"),
   826 => (x"87",x"d4",x"e8",x"49"),
   827 => (x"4c",x"70",x"86",x"c8"),
   828 => (x"06",x"ac",x"b7",x"c0"),
   829 => (x"74",x"87",x"d3",x"c1"),
   830 => (x"49",x"e0",x"c0",x"85"),
   831 => (x"4b",x"75",x"89",x"74"),
   832 => (x"4a",x"c1",x"f8",x"c0"),
   833 => (x"e0",x"cd",x"ff",x"71"),
   834 => (x"c0",x"85",x"c2",x"87"),
   835 => (x"c1",x"48",x"66",x"e4"),
   836 => (x"a6",x"e8",x"c0",x"80"),
   837 => (x"66",x"ec",x"c0",x"58"),
   838 => (x"70",x"81",x"c1",x"49"),
   839 => (x"c8",x"c0",x"02",x"a9"),
   840 => (x"48",x"a6",x"d8",x"87"),
   841 => (x"c5",x"c0",x"78",x"c0"),
   842 => (x"48",x"a6",x"d8",x"87"),
   843 => (x"66",x"d8",x"78",x"c1"),
   844 => (x"49",x"a4",x"c2",x"1e"),
   845 => (x"71",x"48",x"e0",x"c0"),
   846 => (x"1e",x"49",x"70",x"88"),
   847 => (x"ff",x"e6",x"49",x"75"),
   848 => (x"c0",x"86",x"c8",x"87"),
   849 => (x"ff",x"01",x"a8",x"b7"),
   850 => (x"e4",x"c0",x"87",x"c1"),
   851 => (x"d1",x"c0",x"02",x"66"),
   852 => (x"c9",x"49",x"6e",x"87"),
   853 => (x"66",x"e4",x"c0",x"81"),
   854 => (x"c0",x"48",x"6e",x"51"),
   855 => (x"c0",x"78",x"e4",x"e3"),
   856 => (x"49",x"6e",x"87",x"cc"),
   857 => (x"51",x"c2",x"81",x"c9"),
   858 => (x"e4",x"c0",x"48",x"6e"),
   859 => (x"7e",x"c1",x"78",x"d8"),
   860 => (x"e5",x"87",x"c5",x"c0"),
   861 => (x"4c",x"70",x"87",x"f6"),
   862 => (x"f4",x"c0",x"02",x"6e"),
   863 => (x"48",x"66",x"c4",x"87"),
   864 => (x"04",x"a8",x"66",x"c8"),
   865 => (x"c4",x"87",x"cb",x"c0"),
   866 => (x"80",x"c1",x"48",x"66"),
   867 => (x"c0",x"58",x"a6",x"c8"),
   868 => (x"66",x"c8",x"87",x"df"),
   869 => (x"cc",x"88",x"c1",x"48"),
   870 => (x"d4",x"c0",x"58",x"a6"),
   871 => (x"ac",x"c6",x"c1",x"87"),
   872 => (x"87",x"c8",x"c0",x"05"),
   873 => (x"c1",x"48",x"66",x"cc"),
   874 => (x"58",x"a6",x"d0",x"80"),
   875 => (x"70",x"87",x"fd",x"e4"),
   876 => (x"48",x"66",x"d0",x"4c"),
   877 => (x"a6",x"d4",x"80",x"c1"),
   878 => (x"02",x"9c",x"74",x"58"),
   879 => (x"c4",x"87",x"cb",x"c0"),
   880 => (x"c8",x"c1",x"48",x"66"),
   881 => (x"f3",x"04",x"a8",x"66"),
   882 => (x"d6",x"e4",x"87",x"d6"),
   883 => (x"48",x"66",x"c4",x"87"),
   884 => (x"c0",x"03",x"a8",x"c7"),
   885 => (x"f7",x"c1",x"87",x"e5"),
   886 => (x"78",x"c0",x"48",x"c2"),
   887 => (x"cb",x"49",x"66",x"c4"),
   888 => (x"66",x"c0",x"c1",x"91"),
   889 => (x"4a",x"a1",x"c4",x"81"),
   890 => (x"52",x"c0",x"4a",x"6a"),
   891 => (x"48",x"66",x"c4",x"79"),
   892 => (x"a6",x"c8",x"80",x"c1"),
   893 => (x"04",x"a8",x"c7",x"58"),
   894 => (x"ff",x"87",x"db",x"ff"),
   895 => (x"c3",x"ea",x"8e",x"d0"),
   896 => (x"00",x"20",x"3a",x"87"),
   897 => (x"71",x"1e",x"73",x"1e"),
   898 => (x"c6",x"02",x"9b",x"4b"),
   899 => (x"fe",x"f6",x"c1",x"87"),
   900 => (x"c7",x"78",x"c0",x"48"),
   901 => (x"fe",x"f6",x"c1",x"1e"),
   902 => (x"c0",x"1e",x"49",x"bf"),
   903 => (x"c1",x"1e",x"fc",x"f9"),
   904 => (x"49",x"bf",x"fa",x"f6"),
   905 => (x"cc",x"87",x"cc",x"ef"),
   906 => (x"fa",x"f6",x"c1",x"86"),
   907 => (x"cb",x"ea",x"49",x"bf"),
   908 => (x"02",x"9b",x"73",x"87"),
   909 => (x"f9",x"c0",x"87",x"c8"),
   910 => (x"e3",x"c0",x"49",x"fc"),
   911 => (x"c7",x"e9",x"87",x"cb"),
   912 => (x"f9",x"c5",x"1e",x"87"),
   913 => (x"fe",x"49",x"c1",x"87"),
   914 => (x"f0",x"c2",x"87",x"fa"),
   915 => (x"1e",x"4f",x"26",x"87"),
   916 => (x"87",x"d1",x"e7",x"c0"),
   917 => (x"4f",x"26",x"87",x"fa"),
   918 => (x"fe",x"f6",x"c1",x"1e"),
   919 => (x"c1",x"78",x"c0",x"48"),
   920 => (x"c0",x"48",x"fa",x"f6"),
   921 => (x"87",x"d9",x"ff",x"78"),
   922 => (x"48",x"c0",x"87",x"e5"),
   923 => (x"20",x"80",x"4f",x"26"),
   924 => (x"74",x"69",x"78",x"45"),
   925 => (x"42",x"20",x"80",x"00"),
   926 => (x"00",x"6b",x"63",x"61"),
   927 => (x"00",x"00",x"08",x"94"),
   928 => (x"00",x"00",x"1d",x"c6"),
   929 => (x"94",x"00",x"00",x"00"),
   930 => (x"e4",x"00",x"00",x"08"),
   931 => (x"00",x"00",x"00",x"1d"),
   932 => (x"08",x"94",x"00",x"00"),
   933 => (x"1e",x"02",x"00",x"00"),
   934 => (x"00",x"00",x"00",x"00"),
   935 => (x"00",x"08",x"94",x"00"),
   936 => (x"00",x"1e",x"20",x"00"),
   937 => (x"00",x"00",x"00",x"00"),
   938 => (x"00",x"00",x"08",x"94"),
   939 => (x"00",x"00",x"1e",x"3e"),
   940 => (x"94",x"00",x"00",x"00"),
   941 => (x"5c",x"00",x"00",x"08"),
   942 => (x"00",x"00",x"00",x"1e"),
   943 => (x"08",x"94",x"00",x"00"),
   944 => (x"1e",x"7a",x"00",x"00"),
   945 => (x"00",x"00",x"00",x"00"),
   946 => (x"00",x"08",x"94",x"00"),
   947 => (x"00",x"00",x"00",x"00"),
   948 => (x"00",x"00",x"00",x"00"),
   949 => (x"00",x"00",x"09",x"2f"),
   950 => (x"00",x"00",x"00",x"00"),
   951 => (x"4c",x"00",x"00",x"00"),
   952 => (x"20",x"64",x"61",x"6f"),
   953 => (x"1e",x"00",x"2e",x"2a"),
   954 => (x"c0",x"48",x"f0",x"fe"),
   955 => (x"79",x"09",x"cd",x"78"),
   956 => (x"1e",x"4f",x"26",x"09"),
   957 => (x"bf",x"f0",x"fe",x"1e"),
   958 => (x"26",x"26",x"48",x"7e"),
   959 => (x"f0",x"fe",x"1e",x"4f"),
   960 => (x"26",x"78",x"c1",x"48"),
   961 => (x"f0",x"fe",x"1e",x"4f"),
   962 => (x"26",x"78",x"c0",x"48"),
   963 => (x"4a",x"71",x"1e",x"4f"),
   964 => (x"26",x"52",x"52",x"c0"),
   965 => (x"5b",x"5e",x"0e",x"4f"),
   966 => (x"f4",x"0e",x"5d",x"5c"),
   967 => (x"97",x"4d",x"71",x"86"),
   968 => (x"a5",x"c1",x"7e",x"6d"),
   969 => (x"48",x"6c",x"97",x"4c"),
   970 => (x"6e",x"58",x"a6",x"c8"),
   971 => (x"a8",x"66",x"c4",x"48"),
   972 => (x"ff",x"87",x"c5",x"05"),
   973 => (x"87",x"e6",x"c0",x"48"),
   974 => (x"c2",x"87",x"ca",x"ff"),
   975 => (x"6c",x"97",x"49",x"a5"),
   976 => (x"4b",x"a3",x"71",x"4b"),
   977 => (x"97",x"4b",x"6b",x"97"),
   978 => (x"48",x"6e",x"7e",x"6c"),
   979 => (x"a6",x"c8",x"80",x"c1"),
   980 => (x"cc",x"98",x"c7",x"58"),
   981 => (x"97",x"70",x"58",x"a6"),
   982 => (x"87",x"e1",x"fe",x"7c"),
   983 => (x"8e",x"f4",x"48",x"73"),
   984 => (x"4c",x"26",x"4d",x"26"),
   985 => (x"4f",x"26",x"4b",x"26"),
   986 => (x"5c",x"5b",x"5e",x"0e"),
   987 => (x"71",x"86",x"f4",x"0e"),
   988 => (x"4a",x"66",x"d8",x"4c"),
   989 => (x"c2",x"9a",x"ff",x"c3"),
   990 => (x"6c",x"97",x"4b",x"a4"),
   991 => (x"49",x"a1",x"73",x"49"),
   992 => (x"6c",x"97",x"51",x"72"),
   993 => (x"c1",x"48",x"6e",x"7e"),
   994 => (x"58",x"a6",x"c8",x"80"),
   995 => (x"a6",x"cc",x"98",x"c7"),
   996 => (x"f4",x"54",x"70",x"58"),
   997 => (x"87",x"ca",x"ff",x"8e"),
   998 => (x"e8",x"fd",x"1e",x"1e"),
   999 => (x"4a",x"bf",x"e0",x"87"),
  1000 => (x"c0",x"e0",x"c0",x"49"),
  1001 => (x"87",x"cb",x"02",x"99"),
  1002 => (x"fa",x"c1",x"1e",x"72"),
  1003 => (x"f7",x"fe",x"49",x"d8"),
  1004 => (x"fc",x"86",x"c4",x"87"),
  1005 => (x"7e",x"70",x"87",x"fd"),
  1006 => (x"26",x"87",x"c2",x"fd"),
  1007 => (x"c1",x"1e",x"4f",x"26"),
  1008 => (x"fd",x"49",x"d8",x"fa"),
  1009 => (x"fe",x"c0",x"87",x"c7"),
  1010 => (x"da",x"fc",x"49",x"d8"),
  1011 => (x"87",x"d9",x"c5",x"87"),
  1012 => (x"5e",x"0e",x"4f",x"26"),
  1013 => (x"0e",x"5d",x"5c",x"5b"),
  1014 => (x"bf",x"f7",x"fa",x"c1"),
  1015 => (x"e6",x"c0",x"c1",x"4a"),
  1016 => (x"72",x"4c",x"49",x"bf"),
  1017 => (x"fc",x"4d",x"71",x"bc"),
  1018 => (x"4b",x"c0",x"87",x"db"),
  1019 => (x"99",x"d0",x"49",x"74"),
  1020 => (x"75",x"87",x"d5",x"02"),
  1021 => (x"71",x"99",x"d0",x"49"),
  1022 => (x"c1",x"1e",x"c0",x"1e"),
  1023 => (x"73",x"4a",x"f8",x"c6"),
  1024 => (x"c0",x"49",x"12",x"82"),
  1025 => (x"86",x"c8",x"87",x"e4"),
  1026 => (x"83",x"2d",x"2c",x"c1"),
  1027 => (x"ff",x"04",x"ab",x"c8"),
  1028 => (x"e8",x"fb",x"87",x"da"),
  1029 => (x"e6",x"c0",x"c1",x"87"),
  1030 => (x"f7",x"fa",x"c1",x"48"),
  1031 => (x"4d",x"26",x"78",x"bf"),
  1032 => (x"4b",x"26",x"4c",x"26"),
  1033 => (x"00",x"00",x"4f",x"26"),
  1034 => (x"ff",x"1e",x"00",x"00"),
  1035 => (x"e1",x"c8",x"48",x"d0"),
  1036 => (x"48",x"d4",x"ff",x"78"),
  1037 => (x"66",x"c4",x"78",x"c5"),
  1038 => (x"c3",x"87",x"c3",x"02"),
  1039 => (x"66",x"c8",x"78",x"e0"),
  1040 => (x"ff",x"87",x"c6",x"02"),
  1041 => (x"f0",x"c3",x"48",x"d4"),
  1042 => (x"48",x"d4",x"ff",x"78"),
  1043 => (x"d0",x"ff",x"78",x"71"),
  1044 => (x"78",x"e1",x"c8",x"48"),
  1045 => (x"26",x"78",x"e0",x"c0"),
  1046 => (x"5b",x"5e",x"0e",x"4f"),
  1047 => (x"4c",x"71",x"0e",x"5c"),
  1048 => (x"49",x"d8",x"fa",x"c1"),
  1049 => (x"70",x"87",x"ee",x"fa"),
  1050 => (x"aa",x"b7",x"c0",x"4a"),
  1051 => (x"87",x"e3",x"c2",x"04"),
  1052 => (x"05",x"aa",x"e0",x"c3"),
  1053 => (x"c4",x"c1",x"87",x"c9"),
  1054 => (x"78",x"c1",x"48",x"dc"),
  1055 => (x"c3",x"87",x"d4",x"c2"),
  1056 => (x"c9",x"05",x"aa",x"f0"),
  1057 => (x"d8",x"c4",x"c1",x"87"),
  1058 => (x"c1",x"78",x"c1",x"48"),
  1059 => (x"c4",x"c1",x"87",x"f5"),
  1060 => (x"c7",x"02",x"bf",x"dc"),
  1061 => (x"c2",x"4b",x"72",x"87"),
  1062 => (x"87",x"c2",x"b3",x"c0"),
  1063 => (x"9c",x"74",x"4b",x"72"),
  1064 => (x"c1",x"87",x"d1",x"05"),
  1065 => (x"1e",x"bf",x"d8",x"c4"),
  1066 => (x"bf",x"dc",x"c4",x"c1"),
  1067 => (x"fd",x"49",x"72",x"1e"),
  1068 => (x"86",x"c8",x"87",x"f8"),
  1069 => (x"bf",x"d8",x"c4",x"c1"),
  1070 => (x"87",x"e0",x"c0",x"02"),
  1071 => (x"b7",x"c4",x"49",x"73"),
  1072 => (x"c5",x"c1",x"91",x"29"),
  1073 => (x"4a",x"73",x"81",x"f8"),
  1074 => (x"92",x"c2",x"9a",x"cf"),
  1075 => (x"30",x"72",x"48",x"c1"),
  1076 => (x"ba",x"ff",x"4a",x"70"),
  1077 => (x"98",x"69",x"48",x"72"),
  1078 => (x"87",x"db",x"79",x"70"),
  1079 => (x"b7",x"c4",x"49",x"73"),
  1080 => (x"c5",x"c1",x"91",x"29"),
  1081 => (x"4a",x"73",x"81",x"f8"),
  1082 => (x"92",x"c2",x"9a",x"cf"),
  1083 => (x"30",x"72",x"48",x"c3"),
  1084 => (x"69",x"48",x"4a",x"70"),
  1085 => (x"c1",x"79",x"70",x"b0"),
  1086 => (x"c0",x"48",x"dc",x"c4"),
  1087 => (x"d8",x"c4",x"c1",x"78"),
  1088 => (x"c1",x"78",x"c0",x"48"),
  1089 => (x"f8",x"49",x"d8",x"fa"),
  1090 => (x"4a",x"70",x"87",x"cb"),
  1091 => (x"03",x"aa",x"b7",x"c0"),
  1092 => (x"c0",x"87",x"dd",x"fd"),
  1093 => (x"87",x"c8",x"fc",x"48"),
  1094 => (x"00",x"00",x"00",x"00"),
  1095 => (x"00",x"00",x"00",x"00"),
  1096 => (x"49",x"4a",x"71",x"1e"),
  1097 => (x"26",x"87",x"f2",x"fc"),
  1098 => (x"4a",x"c0",x"1e",x"4f"),
  1099 => (x"91",x"c4",x"49",x"72"),
  1100 => (x"81",x"f8",x"c5",x"c1"),
  1101 => (x"82",x"c1",x"79",x"c0"),
  1102 => (x"04",x"aa",x"b7",x"d0"),
  1103 => (x"4f",x"26",x"87",x"ee"),
  1104 => (x"5c",x"5b",x"5e",x"0e"),
  1105 => (x"4d",x"71",x"0e",x"5d"),
  1106 => (x"75",x"87",x"fa",x"f6"),
  1107 => (x"2a",x"b7",x"c4",x"4a"),
  1108 => (x"f8",x"c5",x"c1",x"92"),
  1109 => (x"cf",x"4c",x"75",x"82"),
  1110 => (x"6a",x"94",x"c2",x"9c"),
  1111 => (x"2b",x"74",x"4b",x"49"),
  1112 => (x"48",x"c2",x"9b",x"c3"),
  1113 => (x"4c",x"70",x"30",x"74"),
  1114 => (x"48",x"74",x"bc",x"ff"),
  1115 => (x"7a",x"70",x"98",x"71"),
  1116 => (x"73",x"87",x"ca",x"f6"),
  1117 => (x"87",x"e6",x"fa",x"48"),
  1118 => (x"00",x"00",x"00",x"00"),
  1119 => (x"00",x"00",x"00",x"00"),
  1120 => (x"00",x"00",x"00",x"00"),
  1121 => (x"00",x"00",x"00",x"00"),
  1122 => (x"00",x"00",x"00",x"00"),
  1123 => (x"00",x"00",x"00",x"00"),
  1124 => (x"00",x"00",x"00",x"00"),
  1125 => (x"00",x"00",x"00",x"00"),
  1126 => (x"00",x"00",x"00",x"00"),
  1127 => (x"00",x"00",x"00",x"00"),
  1128 => (x"00",x"00",x"00",x"00"),
  1129 => (x"00",x"00",x"00",x"00"),
  1130 => (x"00",x"00",x"00",x"00"),
  1131 => (x"00",x"00",x"00",x"00"),
  1132 => (x"00",x"00",x"00",x"00"),
  1133 => (x"00",x"00",x"00",x"00"),
  1134 => (x"25",x"26",x"1e",x"16"),
  1135 => (x"3e",x"3d",x"36",x"2e"),
  1136 => (x"48",x"d0",x"ff",x"1e"),
  1137 => (x"71",x"78",x"e1",x"c8"),
  1138 => (x"08",x"d4",x"ff",x"48"),
  1139 => (x"48",x"66",x"c4",x"78"),
  1140 => (x"78",x"08",x"d4",x"ff"),
  1141 => (x"71",x"1e",x"4f",x"26"),
  1142 => (x"1e",x"66",x"c4",x"4a"),
  1143 => (x"49",x"a2",x"e0",x"c1"),
  1144 => (x"c8",x"87",x"dd",x"ff"),
  1145 => (x"b7",x"c8",x"49",x"66"),
  1146 => (x"48",x"d4",x"ff",x"29"),
  1147 => (x"d0",x"ff",x"78",x"71"),
  1148 => (x"78",x"e0",x"c0",x"48"),
  1149 => (x"1e",x"4f",x"26",x"26"),
  1150 => (x"c3",x"4a",x"d4",x"ff"),
  1151 => (x"d0",x"ff",x"7a",x"ff"),
  1152 => (x"78",x"e1",x"c8",x"48"),
  1153 => (x"fa",x"c1",x"7a",x"de"),
  1154 => (x"49",x"7a",x"bf",x"e2"),
  1155 => (x"70",x"28",x"c8",x"48"),
  1156 => (x"d0",x"48",x"71",x"7a"),
  1157 => (x"71",x"7a",x"70",x"28"),
  1158 => (x"70",x"28",x"d8",x"48"),
  1159 => (x"48",x"d0",x"ff",x"7a"),
  1160 => (x"26",x"78",x"e0",x"c0"),
  1161 => (x"5b",x"5e",x"0e",x"4f"),
  1162 => (x"71",x"0e",x"5d",x"5c"),
  1163 => (x"e2",x"fa",x"c1",x"4c"),
  1164 => (x"74",x"4b",x"4d",x"bf"),
  1165 => (x"9b",x"66",x"d0",x"2b"),
  1166 => (x"66",x"d4",x"83",x"c1"),
  1167 => (x"87",x"c2",x"04",x"ab"),
  1168 => (x"4a",x"74",x"4b",x"c0"),
  1169 => (x"72",x"49",x"66",x"d0"),
  1170 => (x"75",x"b9",x"ff",x"31"),
  1171 => (x"72",x"48",x"73",x"99"),
  1172 => (x"48",x"4a",x"70",x"30"),
  1173 => (x"fa",x"c1",x"b0",x"71"),
  1174 => (x"da",x"fe",x"58",x"e6"),
  1175 => (x"26",x"4d",x"26",x"87"),
  1176 => (x"26",x"4b",x"26",x"4c"),
  1177 => (x"d0",x"ff",x"1e",x"4f"),
  1178 => (x"78",x"c9",x"c8",x"48"),
  1179 => (x"d4",x"ff",x"48",x"71"),
  1180 => (x"4f",x"26",x"78",x"08"),
  1181 => (x"49",x"4a",x"71",x"1e"),
  1182 => (x"d0",x"ff",x"87",x"eb"),
  1183 => (x"26",x"78",x"c8",x"48"),
  1184 => (x"1e",x"73",x"1e",x"4f"),
  1185 => (x"fa",x"c1",x"4b",x"71"),
  1186 => (x"c3",x"02",x"bf",x"f2"),
  1187 => (x"87",x"eb",x"c2",x"87"),
  1188 => (x"c8",x"48",x"d0",x"ff"),
  1189 => (x"49",x"73",x"78",x"c9"),
  1190 => (x"ff",x"b1",x"e0",x"c0"),
  1191 => (x"78",x"71",x"48",x"d4"),
  1192 => (x"48",x"e6",x"fa",x"c1"),
  1193 => (x"66",x"c8",x"78",x"c0"),
  1194 => (x"c3",x"87",x"c5",x"02"),
  1195 => (x"87",x"c2",x"49",x"ff"),
  1196 => (x"fa",x"c1",x"49",x"c0"),
  1197 => (x"66",x"cc",x"59",x"ee"),
  1198 => (x"c5",x"87",x"c6",x"02"),
  1199 => (x"c4",x"4a",x"d5",x"d5"),
  1200 => (x"ff",x"ff",x"cf",x"87"),
  1201 => (x"f2",x"fa",x"c1",x"4a"),
  1202 => (x"f2",x"fa",x"c1",x"5a"),
  1203 => (x"c4",x"78",x"c1",x"48"),
  1204 => (x"26",x"4d",x"26",x"87"),
  1205 => (x"26",x"4b",x"26",x"4c"),
  1206 => (x"5b",x"5e",x"0e",x"4f"),
  1207 => (x"71",x"0e",x"5d",x"5c"),
  1208 => (x"ee",x"fa",x"c1",x"4a"),
  1209 => (x"9a",x"72",x"4c",x"bf"),
  1210 => (x"49",x"87",x"cb",x"02"),
  1211 => (x"c9",x"c1",x"91",x"c8"),
  1212 => (x"83",x"71",x"4b",x"f7"),
  1213 => (x"cd",x"c1",x"87",x"c4"),
  1214 => (x"4d",x"c0",x"4b",x"f7"),
  1215 => (x"99",x"74",x"49",x"13"),
  1216 => (x"bf",x"ea",x"fa",x"c1"),
  1217 => (x"48",x"d4",x"ff",x"b9"),
  1218 => (x"b7",x"c1",x"78",x"71"),
  1219 => (x"b7",x"c8",x"85",x"2c"),
  1220 => (x"87",x"e8",x"04",x"ad"),
  1221 => (x"bf",x"e6",x"fa",x"c1"),
  1222 => (x"c1",x"80",x"c8",x"48"),
  1223 => (x"fe",x"58",x"ea",x"fa"),
  1224 => (x"73",x"1e",x"87",x"ef"),
  1225 => (x"13",x"4b",x"71",x"1e"),
  1226 => (x"cb",x"02",x"9a",x"4a"),
  1227 => (x"fe",x"49",x"72",x"87"),
  1228 => (x"4a",x"13",x"87",x"e7"),
  1229 => (x"87",x"f5",x"05",x"9a"),
  1230 => (x"1e",x"87",x"da",x"fe"),
  1231 => (x"bf",x"e6",x"fa",x"c1"),
  1232 => (x"e6",x"fa",x"c1",x"49"),
  1233 => (x"78",x"a1",x"c1",x"48"),
  1234 => (x"a9",x"b7",x"c0",x"c4"),
  1235 => (x"ff",x"87",x"db",x"03"),
  1236 => (x"fa",x"c1",x"48",x"d4"),
  1237 => (x"c1",x"78",x"bf",x"ea"),
  1238 => (x"49",x"bf",x"e6",x"fa"),
  1239 => (x"48",x"e6",x"fa",x"c1"),
  1240 => (x"c4",x"78",x"a1",x"c1"),
  1241 => (x"04",x"a9",x"b7",x"c0"),
  1242 => (x"d0",x"ff",x"87",x"e5"),
  1243 => (x"c1",x"78",x"c8",x"48"),
  1244 => (x"c0",x"48",x"f2",x"fa"),
  1245 => (x"00",x"4f",x"26",x"78"),
  1246 => (x"00",x"00",x"00",x"00"),
  1247 => (x"00",x"00",x"00",x"00"),
  1248 => (x"5f",x"5f",x"00",x"00"),
  1249 => (x"00",x"00",x"00",x"00"),
  1250 => (x"03",x"00",x"03",x"03"),
  1251 => (x"14",x"00",x"00",x"03"),
  1252 => (x"7f",x"14",x"7f",x"7f"),
  1253 => (x"00",x"00",x"14",x"7f"),
  1254 => (x"6b",x"6b",x"2e",x"24"),
  1255 => (x"4c",x"00",x"12",x"3a"),
  1256 => (x"6c",x"18",x"36",x"6a"),
  1257 => (x"30",x"00",x"32",x"56"),
  1258 => (x"77",x"59",x"4f",x"7e"),
  1259 => (x"00",x"40",x"68",x"3a"),
  1260 => (x"03",x"07",x"04",x"00"),
  1261 => (x"00",x"00",x"00",x"00"),
  1262 => (x"63",x"3e",x"1c",x"00"),
  1263 => (x"00",x"00",x"00",x"41"),
  1264 => (x"3e",x"63",x"41",x"00"),
  1265 => (x"08",x"00",x"00",x"1c"),
  1266 => (x"1c",x"1c",x"3e",x"2a"),
  1267 => (x"00",x"08",x"2a",x"3e"),
  1268 => (x"3e",x"3e",x"08",x"08"),
  1269 => (x"00",x"00",x"08",x"08"),
  1270 => (x"60",x"e0",x"80",x"00"),
  1271 => (x"00",x"00",x"00",x"00"),
  1272 => (x"08",x"08",x"08",x"08"),
  1273 => (x"00",x"00",x"08",x"08"),
  1274 => (x"60",x"60",x"00",x"00"),
  1275 => (x"40",x"00",x"00",x"00"),
  1276 => (x"0c",x"18",x"30",x"60"),
  1277 => (x"00",x"01",x"03",x"06"),
  1278 => (x"4d",x"59",x"7f",x"3e"),
  1279 => (x"00",x"00",x"3e",x"7f"),
  1280 => (x"7f",x"7f",x"06",x"04"),
  1281 => (x"00",x"00",x"00",x"00"),
  1282 => (x"59",x"71",x"63",x"42"),
  1283 => (x"00",x"00",x"46",x"4f"),
  1284 => (x"49",x"49",x"63",x"22"),
  1285 => (x"18",x"00",x"36",x"7f"),
  1286 => (x"7f",x"13",x"16",x"1c"),
  1287 => (x"00",x"00",x"10",x"7f"),
  1288 => (x"45",x"45",x"67",x"27"),
  1289 => (x"00",x"00",x"39",x"7d"),
  1290 => (x"49",x"4b",x"7e",x"3c"),
  1291 => (x"00",x"00",x"30",x"79"),
  1292 => (x"79",x"71",x"01",x"01"),
  1293 => (x"00",x"00",x"07",x"0f"),
  1294 => (x"49",x"49",x"7f",x"36"),
  1295 => (x"00",x"00",x"36",x"7f"),
  1296 => (x"69",x"49",x"4f",x"06"),
  1297 => (x"00",x"00",x"1e",x"3f"),
  1298 => (x"66",x"66",x"00",x"00"),
  1299 => (x"00",x"00",x"00",x"00"),
  1300 => (x"66",x"e6",x"80",x"00"),
  1301 => (x"00",x"00",x"00",x"00"),
  1302 => (x"14",x"14",x"08",x"08"),
  1303 => (x"00",x"00",x"22",x"22"),
  1304 => (x"14",x"14",x"14",x"14"),
  1305 => (x"00",x"00",x"14",x"14"),
  1306 => (x"14",x"14",x"22",x"22"),
  1307 => (x"00",x"00",x"08",x"08"),
  1308 => (x"59",x"51",x"03",x"02"),
  1309 => (x"3e",x"00",x"06",x"0f"),
  1310 => (x"55",x"5d",x"41",x"7f"),
  1311 => (x"00",x"00",x"1e",x"1f"),
  1312 => (x"09",x"09",x"7f",x"7e"),
  1313 => (x"00",x"00",x"7e",x"7f"),
  1314 => (x"49",x"49",x"7f",x"7f"),
  1315 => (x"00",x"00",x"36",x"7f"),
  1316 => (x"41",x"63",x"3e",x"1c"),
  1317 => (x"00",x"00",x"41",x"41"),
  1318 => (x"63",x"41",x"7f",x"7f"),
  1319 => (x"00",x"00",x"1c",x"3e"),
  1320 => (x"49",x"49",x"7f",x"7f"),
  1321 => (x"00",x"00",x"41",x"41"),
  1322 => (x"09",x"09",x"7f",x"7f"),
  1323 => (x"00",x"00",x"01",x"01"),
  1324 => (x"49",x"41",x"7f",x"3e"),
  1325 => (x"00",x"00",x"7a",x"7b"),
  1326 => (x"08",x"08",x"7f",x"7f"),
  1327 => (x"00",x"00",x"7f",x"7f"),
  1328 => (x"7f",x"7f",x"41",x"00"),
  1329 => (x"00",x"00",x"00",x"41"),
  1330 => (x"40",x"40",x"60",x"20"),
  1331 => (x"7f",x"00",x"3f",x"7f"),
  1332 => (x"36",x"1c",x"08",x"7f"),
  1333 => (x"00",x"00",x"41",x"63"),
  1334 => (x"40",x"40",x"7f",x"7f"),
  1335 => (x"7f",x"00",x"40",x"40"),
  1336 => (x"06",x"0c",x"06",x"7f"),
  1337 => (x"7f",x"00",x"7f",x"7f"),
  1338 => (x"18",x"0c",x"06",x"7f"),
  1339 => (x"00",x"00",x"7f",x"7f"),
  1340 => (x"41",x"41",x"7f",x"3e"),
  1341 => (x"00",x"00",x"3e",x"7f"),
  1342 => (x"09",x"09",x"7f",x"7f"),
  1343 => (x"3e",x"00",x"06",x"0f"),
  1344 => (x"7f",x"61",x"41",x"7f"),
  1345 => (x"00",x"00",x"40",x"7e"),
  1346 => (x"19",x"09",x"7f",x"7f"),
  1347 => (x"00",x"00",x"66",x"7f"),
  1348 => (x"59",x"4d",x"6f",x"26"),
  1349 => (x"00",x"00",x"32",x"7b"),
  1350 => (x"7f",x"7f",x"01",x"01"),
  1351 => (x"00",x"00",x"01",x"01"),
  1352 => (x"40",x"40",x"7f",x"3f"),
  1353 => (x"00",x"00",x"3f",x"7f"),
  1354 => (x"70",x"70",x"3f",x"0f"),
  1355 => (x"7f",x"00",x"0f",x"3f"),
  1356 => (x"30",x"18",x"30",x"7f"),
  1357 => (x"41",x"00",x"7f",x"7f"),
  1358 => (x"1c",x"1c",x"36",x"63"),
  1359 => (x"01",x"41",x"63",x"36"),
  1360 => (x"7c",x"7c",x"06",x"03"),
  1361 => (x"61",x"01",x"03",x"06"),
  1362 => (x"47",x"4d",x"59",x"71"),
  1363 => (x"00",x"00",x"41",x"43"),
  1364 => (x"41",x"7f",x"7f",x"00"),
  1365 => (x"01",x"00",x"00",x"41"),
  1366 => (x"18",x"0c",x"06",x"03"),
  1367 => (x"00",x"40",x"60",x"30"),
  1368 => (x"7f",x"41",x"41",x"00"),
  1369 => (x"08",x"00",x"00",x"7f"),
  1370 => (x"06",x"03",x"06",x"0c"),
  1371 => (x"80",x"00",x"08",x"0c"),
  1372 => (x"80",x"80",x"80",x"80"),
  1373 => (x"00",x"00",x"80",x"80"),
  1374 => (x"07",x"03",x"00",x"00"),
  1375 => (x"00",x"00",x"00",x"04"),
  1376 => (x"54",x"54",x"74",x"20"),
  1377 => (x"00",x"00",x"78",x"7c"),
  1378 => (x"44",x"44",x"7f",x"7f"),
  1379 => (x"00",x"00",x"38",x"7c"),
  1380 => (x"44",x"44",x"7c",x"38"),
  1381 => (x"00",x"00",x"00",x"44"),
  1382 => (x"44",x"44",x"7c",x"38"),
  1383 => (x"00",x"00",x"7f",x"7f"),
  1384 => (x"54",x"54",x"7c",x"38"),
  1385 => (x"00",x"00",x"18",x"5c"),
  1386 => (x"05",x"7f",x"7e",x"04"),
  1387 => (x"00",x"00",x"00",x"05"),
  1388 => (x"a4",x"a4",x"bc",x"18"),
  1389 => (x"00",x"00",x"7c",x"fc"),
  1390 => (x"04",x"04",x"7f",x"7f"),
  1391 => (x"00",x"00",x"78",x"7c"),
  1392 => (x"7d",x"3d",x"00",x"00"),
  1393 => (x"00",x"00",x"00",x"40"),
  1394 => (x"fd",x"80",x"80",x"80"),
  1395 => (x"00",x"00",x"00",x"7d"),
  1396 => (x"38",x"10",x"7f",x"7f"),
  1397 => (x"00",x"00",x"44",x"6c"),
  1398 => (x"7f",x"3f",x"00",x"00"),
  1399 => (x"7c",x"00",x"00",x"40"),
  1400 => (x"0c",x"18",x"0c",x"7c"),
  1401 => (x"00",x"00",x"78",x"7c"),
  1402 => (x"04",x"04",x"7c",x"7c"),
  1403 => (x"00",x"00",x"78",x"7c"),
  1404 => (x"44",x"44",x"7c",x"38"),
  1405 => (x"00",x"00",x"38",x"7c"),
  1406 => (x"24",x"24",x"fc",x"fc"),
  1407 => (x"00",x"00",x"18",x"3c"),
  1408 => (x"24",x"24",x"3c",x"18"),
  1409 => (x"00",x"00",x"fc",x"fc"),
  1410 => (x"04",x"04",x"7c",x"7c"),
  1411 => (x"00",x"00",x"08",x"0c"),
  1412 => (x"54",x"54",x"5c",x"48"),
  1413 => (x"00",x"00",x"20",x"74"),
  1414 => (x"44",x"7f",x"3f",x"04"),
  1415 => (x"00",x"00",x"00",x"44"),
  1416 => (x"40",x"40",x"7c",x"3c"),
  1417 => (x"00",x"00",x"7c",x"7c"),
  1418 => (x"60",x"60",x"3c",x"1c"),
  1419 => (x"3c",x"00",x"1c",x"3c"),
  1420 => (x"60",x"30",x"60",x"7c"),
  1421 => (x"44",x"00",x"3c",x"7c"),
  1422 => (x"38",x"10",x"38",x"6c"),
  1423 => (x"00",x"00",x"44",x"6c"),
  1424 => (x"60",x"e0",x"bc",x"1c"),
  1425 => (x"00",x"00",x"1c",x"3c"),
  1426 => (x"5c",x"74",x"64",x"44"),
  1427 => (x"00",x"00",x"44",x"4c"),
  1428 => (x"77",x"3e",x"08",x"08"),
  1429 => (x"00",x"00",x"41",x"41"),
  1430 => (x"7f",x"7f",x"00",x"00"),
  1431 => (x"00",x"00",x"00",x"00"),
  1432 => (x"3e",x"77",x"41",x"41"),
  1433 => (x"02",x"00",x"08",x"08"),
  1434 => (x"02",x"03",x"01",x"01"),
  1435 => (x"7f",x"00",x"01",x"02"),
  1436 => (x"7f",x"7f",x"7f",x"7f"),
  1437 => (x"08",x"00",x"7f",x"7f"),
  1438 => (x"3e",x"1c",x"1c",x"08"),
  1439 => (x"7f",x"7f",x"7f",x"3e"),
  1440 => (x"1c",x"3e",x"3e",x"7f"),
  1441 => (x"00",x"08",x"08",x"1c"),
  1442 => (x"7c",x"7c",x"18",x"10"),
  1443 => (x"00",x"00",x"10",x"18"),
  1444 => (x"7c",x"7c",x"30",x"10"),
  1445 => (x"10",x"00",x"10",x"30"),
  1446 => (x"78",x"60",x"60",x"30"),
  1447 => (x"42",x"00",x"06",x"1e"),
  1448 => (x"3c",x"18",x"3c",x"66"),
  1449 => (x"78",x"00",x"42",x"66"),
  1450 => (x"c6",x"c2",x"6a",x"38"),
  1451 => (x"60",x"00",x"38",x"6c"),
  1452 => (x"00",x"60",x"00",x"00"),
  1453 => (x"0e",x"00",x"60",x"00"),
  1454 => (x"5d",x"5c",x"5b",x"5e"),
  1455 => (x"4c",x"71",x"1e",x"0e"),
  1456 => (x"bf",x"c3",x"fb",x"c1"),
  1457 => (x"c0",x"4b",x"c0",x"4d"),
  1458 => (x"02",x"ab",x"74",x"1e"),
  1459 => (x"a6",x"c4",x"87",x"c7"),
  1460 => (x"c5",x"78",x"c0",x"48"),
  1461 => (x"48",x"a6",x"c4",x"87"),
  1462 => (x"66",x"c4",x"78",x"c1"),
  1463 => (x"ee",x"49",x"73",x"1e"),
  1464 => (x"86",x"c8",x"87",x"df"),
  1465 => (x"ef",x"49",x"e0",x"c0"),
  1466 => (x"a5",x"c4",x"87",x"ef"),
  1467 => (x"f0",x"49",x"6a",x"4a"),
  1468 => (x"c6",x"f1",x"87",x"f0"),
  1469 => (x"c1",x"85",x"cb",x"87"),
  1470 => (x"ab",x"b7",x"c8",x"83"),
  1471 => (x"87",x"c7",x"ff",x"04"),
  1472 => (x"26",x"4d",x"26",x"26"),
  1473 => (x"26",x"4b",x"26",x"4c"),
  1474 => (x"4a",x"71",x"1e",x"4f"),
  1475 => (x"5a",x"c7",x"fb",x"c1"),
  1476 => (x"48",x"c7",x"fb",x"c1"),
  1477 => (x"fe",x"49",x"78",x"c7"),
  1478 => (x"4f",x"26",x"87",x"dd"),
  1479 => (x"71",x"1e",x"73",x"1e"),
  1480 => (x"aa",x"b7",x"c0",x"4a"),
  1481 => (x"c1",x"87",x"d3",x"03"),
  1482 => (x"05",x"bf",x"db",x"e8"),
  1483 => (x"4b",x"c1",x"87",x"c4"),
  1484 => (x"4b",x"c0",x"87",x"c2"),
  1485 => (x"5b",x"df",x"e8",x"c1"),
  1486 => (x"e8",x"c1",x"87",x"c4"),
  1487 => (x"e8",x"c1",x"5a",x"df"),
  1488 => (x"c1",x"4a",x"bf",x"db"),
  1489 => (x"a2",x"c0",x"c1",x"9a"),
  1490 => (x"87",x"e8",x"ec",x"49"),
  1491 => (x"e8",x"c1",x"48",x"fc"),
  1492 => (x"fe",x"78",x"bf",x"db"),
  1493 => (x"71",x"1e",x"87",x"ef"),
  1494 => (x"1e",x"66",x"c4",x"4a"),
  1495 => (x"f5",x"e9",x"49",x"72"),
  1496 => (x"4f",x"26",x"26",x"87"),
  1497 => (x"db",x"e8",x"c1",x"1e"),
  1498 => (x"f3",x"e6",x"49",x"bf"),
  1499 => (x"fb",x"fa",x"c1",x"87"),
  1500 => (x"78",x"bf",x"e8",x"48"),
  1501 => (x"48",x"f7",x"fa",x"c1"),
  1502 => (x"c1",x"78",x"bf",x"ec"),
  1503 => (x"4a",x"bf",x"fb",x"fa"),
  1504 => (x"99",x"ff",x"c3",x"49"),
  1505 => (x"72",x"2a",x"b7",x"c8"),
  1506 => (x"c1",x"b0",x"71",x"48"),
  1507 => (x"26",x"58",x"c3",x"fb"),
  1508 => (x"5b",x"5e",x"0e",x"4f"),
  1509 => (x"71",x"0e",x"5d",x"5c"),
  1510 => (x"87",x"c8",x"ff",x"4b"),
  1511 => (x"48",x"f6",x"fa",x"c1"),
  1512 => (x"49",x"73",x"50",x"c0"),
  1513 => (x"70",x"87",x"d9",x"e6"),
  1514 => (x"9c",x"c2",x"4c",x"49"),
  1515 => (x"c9",x"49",x"ee",x"cb"),
  1516 => (x"49",x"70",x"87",x"f1"),
  1517 => (x"f6",x"fa",x"c1",x"4d"),
  1518 => (x"c1",x"05",x"bf",x"97"),
  1519 => (x"66",x"d0",x"87",x"e2"),
  1520 => (x"ff",x"fa",x"c1",x"49"),
  1521 => (x"d6",x"05",x"99",x"bf"),
  1522 => (x"49",x"66",x"d4",x"87"),
  1523 => (x"bf",x"f7",x"fa",x"c1"),
  1524 => (x"87",x"cb",x"05",x"99"),
  1525 => (x"e7",x"e5",x"49",x"73"),
  1526 => (x"02",x"98",x"70",x"87"),
  1527 => (x"c1",x"87",x"c1",x"c1"),
  1528 => (x"87",x"c0",x"fe",x"4c"),
  1529 => (x"c6",x"c9",x"49",x"75"),
  1530 => (x"02",x"98",x"70",x"87"),
  1531 => (x"fa",x"c1",x"87",x"c6"),
  1532 => (x"50",x"c1",x"48",x"f6"),
  1533 => (x"97",x"f6",x"fa",x"c1"),
  1534 => (x"e3",x"c0",x"05",x"bf"),
  1535 => (x"ff",x"fa",x"c1",x"87"),
  1536 => (x"66",x"d0",x"49",x"bf"),
  1537 => (x"d6",x"ff",x"05",x"99"),
  1538 => (x"f7",x"fa",x"c1",x"87"),
  1539 => (x"66",x"d4",x"49",x"bf"),
  1540 => (x"ca",x"ff",x"05",x"99"),
  1541 => (x"e4",x"49",x"73",x"87"),
  1542 => (x"98",x"70",x"87",x"e6"),
  1543 => (x"87",x"ff",x"fe",x"05"),
  1544 => (x"dc",x"fb",x"48",x"74"),
  1545 => (x"5b",x"5e",x"0e",x"87"),
  1546 => (x"f4",x"0e",x"5d",x"5c"),
  1547 => (x"4c",x"4d",x"c0",x"86"),
  1548 => (x"c4",x"7e",x"bf",x"ec"),
  1549 => (x"fb",x"c1",x"48",x"a6"),
  1550 => (x"c1",x"78",x"bf",x"c3"),
  1551 => (x"c7",x"1e",x"c0",x"1e"),
  1552 => (x"87",x"cd",x"fd",x"49"),
  1553 => (x"98",x"70",x"86",x"c8"),
  1554 => (x"ff",x"87",x"cd",x"02"),
  1555 => (x"87",x"cc",x"fb",x"49"),
  1556 => (x"e3",x"49",x"da",x"c1"),
  1557 => (x"4d",x"c1",x"87",x"ea"),
  1558 => (x"97",x"f6",x"fa",x"c1"),
  1559 => (x"87",x"c3",x"02",x"bf"),
  1560 => (x"c1",x"87",x"e5",x"c7"),
  1561 => (x"4b",x"bf",x"fb",x"fa"),
  1562 => (x"bf",x"db",x"e8",x"c1"),
  1563 => (x"87",x"e9",x"c0",x"05"),
  1564 => (x"e3",x"49",x"fd",x"c3"),
  1565 => (x"fa",x"c3",x"87",x"ca"),
  1566 => (x"87",x"c4",x"e3",x"49"),
  1567 => (x"ff",x"c3",x"49",x"73"),
  1568 => (x"c0",x"1e",x"71",x"99"),
  1569 => (x"87",x"ce",x"fb",x"49"),
  1570 => (x"b7",x"c8",x"49",x"73"),
  1571 => (x"c1",x"1e",x"71",x"29"),
  1572 => (x"87",x"c2",x"fb",x"49"),
  1573 => (x"f9",x"c5",x"86",x"c8"),
  1574 => (x"ff",x"fa",x"c1",x"87"),
  1575 => (x"02",x"9b",x"4b",x"bf"),
  1576 => (x"e8",x"c1",x"87",x"dd"),
  1577 => (x"c6",x"49",x"bf",x"d7"),
  1578 => (x"98",x"70",x"87",x"c5"),
  1579 => (x"c0",x"87",x"c4",x"05"),
  1580 => (x"c2",x"87",x"d2",x"4b"),
  1581 => (x"ea",x"c5",x"49",x"e0"),
  1582 => (x"db",x"e8",x"c1",x"87"),
  1583 => (x"c1",x"87",x"c6",x"58"),
  1584 => (x"c0",x"48",x"d7",x"e8"),
  1585 => (x"c2",x"49",x"73",x"78"),
  1586 => (x"87",x"cd",x"05",x"99"),
  1587 => (x"e1",x"49",x"eb",x"c3"),
  1588 => (x"49",x"70",x"87",x"ee"),
  1589 => (x"c2",x"02",x"99",x"c2"),
  1590 => (x"73",x"4c",x"fb",x"87"),
  1591 => (x"05",x"99",x"c1",x"49"),
  1592 => (x"f4",x"c3",x"87",x"cd"),
  1593 => (x"87",x"d8",x"e1",x"49"),
  1594 => (x"99",x"c2",x"49",x"70"),
  1595 => (x"fa",x"87",x"c2",x"02"),
  1596 => (x"c8",x"49",x"73",x"4c"),
  1597 => (x"87",x"cd",x"05",x"99"),
  1598 => (x"e1",x"49",x"f5",x"c3"),
  1599 => (x"49",x"70",x"87",x"c2"),
  1600 => (x"d4",x"02",x"99",x"c2"),
  1601 => (x"c7",x"fb",x"c1",x"87"),
  1602 => (x"87",x"c9",x"02",x"bf"),
  1603 => (x"c1",x"88",x"c1",x"48"),
  1604 => (x"c2",x"58",x"cb",x"fb"),
  1605 => (x"c1",x"4c",x"ff",x"87"),
  1606 => (x"c4",x"49",x"73",x"4d"),
  1607 => (x"87",x"cd",x"05",x"99"),
  1608 => (x"e0",x"49",x"f2",x"c3"),
  1609 => (x"49",x"70",x"87",x"da"),
  1610 => (x"db",x"02",x"99",x"c2"),
  1611 => (x"c7",x"fb",x"c1",x"87"),
  1612 => (x"c7",x"48",x"7e",x"bf"),
  1613 => (x"cb",x"03",x"a8",x"b7"),
  1614 => (x"c1",x"48",x"6e",x"87"),
  1615 => (x"cb",x"fb",x"c1",x"80"),
  1616 => (x"87",x"c2",x"c0",x"58"),
  1617 => (x"4d",x"c1",x"4c",x"fe"),
  1618 => (x"ff",x"49",x"fd",x"c3"),
  1619 => (x"70",x"87",x"f1",x"df"),
  1620 => (x"02",x"99",x"c2",x"49"),
  1621 => (x"fb",x"c1",x"87",x"d5"),
  1622 => (x"c0",x"02",x"bf",x"c7"),
  1623 => (x"fb",x"c1",x"87",x"c9"),
  1624 => (x"78",x"c0",x"48",x"c7"),
  1625 => (x"fd",x"87",x"c2",x"c0"),
  1626 => (x"c3",x"4d",x"c1",x"4c"),
  1627 => (x"df",x"ff",x"49",x"fa"),
  1628 => (x"49",x"70",x"87",x"ce"),
  1629 => (x"d9",x"02",x"99",x"c2"),
  1630 => (x"c7",x"fb",x"c1",x"87"),
  1631 => (x"b7",x"c7",x"48",x"bf"),
  1632 => (x"c9",x"c0",x"03",x"a8"),
  1633 => (x"c7",x"fb",x"c1",x"87"),
  1634 => (x"c0",x"78",x"c7",x"48"),
  1635 => (x"4c",x"fc",x"87",x"c2"),
  1636 => (x"b7",x"c0",x"4d",x"c1"),
  1637 => (x"d1",x"c0",x"03",x"ac"),
  1638 => (x"4a",x"66",x"c4",x"87"),
  1639 => (x"6a",x"82",x"d8",x"c1"),
  1640 => (x"87",x"c6",x"c0",x"02"),
  1641 => (x"49",x"74",x"4b",x"6a"),
  1642 => (x"1e",x"c0",x"0f",x"73"),
  1643 => (x"c1",x"1e",x"f0",x"c3"),
  1644 => (x"dc",x"f7",x"49",x"da"),
  1645 => (x"70",x"86",x"c8",x"87"),
  1646 => (x"e2",x"c0",x"02",x"98"),
  1647 => (x"48",x"a6",x"c8",x"87"),
  1648 => (x"bf",x"c7",x"fb",x"c1"),
  1649 => (x"49",x"66",x"c8",x"78"),
  1650 => (x"66",x"c4",x"91",x"cb"),
  1651 => (x"70",x"80",x"71",x"48"),
  1652 => (x"02",x"bf",x"6e",x"7e"),
  1653 => (x"6e",x"87",x"c8",x"c0"),
  1654 => (x"66",x"c8",x"4b",x"bf"),
  1655 => (x"75",x"0f",x"73",x"49"),
  1656 => (x"c8",x"c0",x"02",x"9d"),
  1657 => (x"c7",x"fb",x"c1",x"87"),
  1658 => (x"ca",x"f3",x"49",x"bf"),
  1659 => (x"df",x"e8",x"c1",x"87"),
  1660 => (x"dd",x"c0",x"02",x"bf"),
  1661 => (x"f6",x"c0",x"49",x"87"),
  1662 => (x"02",x"98",x"70",x"87"),
  1663 => (x"c1",x"87",x"d3",x"c0"),
  1664 => (x"49",x"bf",x"c7",x"fb"),
  1665 => (x"c0",x"87",x"f0",x"f2"),
  1666 => (x"87",x"d0",x"f4",x"49"),
  1667 => (x"48",x"df",x"e8",x"c1"),
  1668 => (x"8e",x"f4",x"78",x"c0"),
  1669 => (x"00",x"87",x"ea",x"f3"),
  1670 => (x"00",x"00",x"00",x"00"),
  1671 => (x"00",x"00",x"00",x"00"),
  1672 => (x"1e",x"00",x"00",x"00"),
  1673 => (x"c8",x"ff",x"4a",x"71"),
  1674 => (x"a1",x"72",x"49",x"bf"),
  1675 => (x"1e",x"4f",x"26",x"48"),
  1676 => (x"89",x"bf",x"c8",x"ff"),
  1677 => (x"c0",x"c0",x"c0",x"fe"),
  1678 => (x"01",x"a9",x"c0",x"c0"),
  1679 => (x"4a",x"c0",x"87",x"c4"),
  1680 => (x"4a",x"c1",x"87",x"c2"),
  1681 => (x"4f",x"26",x"48",x"72"),
  1682 => (x"f1",x"e9",x"c1",x"1e"),
  1683 => (x"b9",x"c1",x"49",x"bf"),
  1684 => (x"59",x"f5",x"e9",x"c1"),
  1685 => (x"c3",x"48",x"d4",x"ff"),
  1686 => (x"d0",x"ff",x"78",x"ff"),
  1687 => (x"78",x"e1",x"c8",x"48"),
  1688 => (x"c1",x"48",x"d4",x"ff"),
  1689 => (x"71",x"31",x"c4",x"78"),
  1690 => (x"48",x"d0",x"ff",x"78"),
  1691 => (x"26",x"78",x"e0",x"c0"),
  1692 => (x"00",x"00",x"00",x"4f"),
  1693 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

